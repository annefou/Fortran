netcdf \2t_20140623 {
dimensions:
	x = 161 ;
	y = 286 ;
variables:
	float T2M(x, y) ;
		T2M:long_name = "2 metre temperature" ;
		T2M:units = "K" ;
		T2M:code = 167 ;
		T2M:table = 128 ;

// global attributes:
		:CDI = "Climate Data Interface version 1.7.0 (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "Mon Mar 14 10:00:04 2016: cdo -t ecmwf -f nc copy 2t_20140623_12.grib 2t_20140623.nc" ;
		:institution = "European Centre for Medium-Range Weather Forecasts" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 T2M =
  274.9001, 274.9072, 274.9141, 274.9209, 274.9277, 274.9348, 274.9417, 
    274.9558, 275.0212, 275.0864, 275.1519, 275.217, 275.2825, 275.3477, 
    275.4131, 275.4785, 275.5437, 275.6091, 275.6743, 275.7397, 275.8049, 
    275.875, 276.0127, 276.1506, 276.2883, 276.4263, 276.5642, 276.7019, 
    276.8398, 276.9775, 277.1155, 277.2534, 277.3911, 277.5291, 277.6667, 
    277.8047, 277.8582, 277.9116, 277.9651, 278.0188, 278.0723, 278.1257, 
    278.1792, 278.2327, 278.2861, 278.3398, 278.3933, 278.4468, 278.5002, 
    278.5537, 278.4966, 278.4319, 278.3672, 278.3025, 278.238, 278.1733, 
    278.1086, 278.0439, 277.9792, 277.9148, 277.8501, 277.7854, 277.7207, 
    277.6562, 277.6853, 277.7278, 277.7703, 277.8127, 277.8552, 277.8977, 
    277.9402, 277.9827, 278.0251, 278.0676, 278.1101, 278.1523, 278.1948, 
    278.2373, 278.3286, 278.4312, 278.5337, 278.636, 278.7385, 278.8411, 
    278.9436, 279.0459, 279.1484, 279.251, 279.3535, 279.4558, 279.5583, 
    279.6609, 279.76, 279.8577, 279.9556, 280.0535, 280.1514, 280.2493, 
    280.3472, 280.4451, 280.543, 280.6409, 280.7388, 280.8367, 280.9346, 
    281.0325, 281.0791, 281.1021, 281.1252, 281.1482, 281.1714, 281.1943, 
    281.2175, 281.2407, 281.2637, 281.2869, 281.3098, 281.333, 281.356, 
    281.3792, 281.3398, 281.2629, 281.186, 281.1091, 281.0325, 280.9556, 
    280.8787, 280.802, 280.7251, 280.6482, 280.5713, 280.4946, 280.4177, 
    280.3408, 280.2922, 280.2659, 280.2393, 280.2126, 280.1863, 280.1597, 
    280.1331, 280.1067, 280.0801, 280.0535, 280.0271, 280.0005, 279.9739, 
    279.9475, 279.9683, 280.0366, 280.1047, 280.1731, 280.2415, 280.3096, 
    280.3779, 280.4463, 280.5144, 280.5828, 280.6509, 280.7192, 280.7876, 
    280.8557, 280.8694, 280.8123, 280.7554, 280.6985, 280.6416, 280.5847, 
    280.5276, 280.4707, 280.4138, 280.3569, 280.3, 280.2432, 280.186, 
    280.1292, 280.0815, 280.0491, 280.0166, 279.9841, 279.9517, 279.9192, 
    279.887, 279.8545, 279.822, 279.7896, 279.7571, 279.7249, 279.6924, 
    279.6599, 279.6497, 279.688, 279.7266, 279.7649, 279.8035, 279.8418, 
    279.8804, 279.9187, 279.9573, 279.9958, 280.0342, 280.0728, 280.1111, 
    280.1497, 280.1697, 280.1348, 280.0999, 280.0647, 280.0298, 279.9949, 
    279.96, 279.925, 279.8899, 279.855, 279.8201, 279.7852, 279.7502, 
    279.7153, 279.6736, 279.6028, 279.532, 279.4612, 279.3906, 279.3198, 
    279.249, 279.1782, 279.1074, 279.0366, 278.9661, 278.8953, 278.8245, 
    278.7537, 278.6885, 278.6614, 278.6343, 278.6072, 278.5801, 278.553, 
    278.5259, 278.4988, 278.4717, 278.4446, 278.4175, 278.3904, 278.3633, 
    278.3362, 278.3113, 278.3181, 278.325, 278.3318, 278.3389, 278.3457, 
    278.3525, 278.3594, 278.3662, 278.3733, 278.3801, 278.387, 278.3938, 
    278.4006, 278.4077, 278.4104, 278.4133, 278.4163, 278.4189, 278.4219, 
    278.4248, 278.4275, 278.4304, 278.4333, 278.436, 278.439, 278.4419, 
    278.4446, 278.4475, 278.4038, 278.3572, 278.3105, 278.2639, 278.217, 
    278.1704, 278.1238, 278.0771, 278.0305, 277.9836, 277.937,
  274.8982, 274.9099, 274.9216, 274.9336, 274.9453, 274.9573, 274.969, 
    274.9863, 275.043, 275.0996, 275.1562, 275.2129, 275.2695, 275.3262, 
    275.3831, 275.4397, 275.4963, 275.553, 275.6096, 275.6663, 275.7229, 
    275.7837, 275.9058, 276.0278, 276.1499, 276.272, 276.394, 276.5161, 
    276.6382, 276.7603, 276.8823, 277.0044, 277.1267, 277.2488, 277.3708, 
    277.4929, 277.5608, 277.6289, 277.697, 277.7649, 277.833, 277.9011, 
    277.969, 278.0371, 278.1052, 278.1731, 278.2412, 278.3093, 278.3772, 
    278.4453, 278.4082, 278.364, 278.3198, 278.2754, 278.2312, 278.187, 
    278.1428, 278.0986, 278.0544, 278.0103, 277.9661, 277.9219, 277.8777, 
    277.8333, 277.864, 277.9053, 277.9465, 277.9878, 278.0291, 278.0703, 
    278.1118, 278.1531, 278.1943, 278.2356, 278.2769, 278.3181, 278.3594, 
    278.4009, 278.4839, 278.5764, 278.6692, 278.7617, 278.8545, 278.9473, 
    279.0398, 279.1326, 279.2251, 279.3179, 279.4106, 279.5032, 279.5959, 
    279.6885, 279.782, 279.8755, 279.969, 280.0625, 280.156, 280.2495, 
    280.343, 280.4365, 280.53, 280.6235, 280.7173, 280.8108, 280.9043, 
    280.9978, 281.0547, 281.095, 281.135, 281.1753, 281.2156, 281.2559, 
    281.2959, 281.3362, 281.3765, 281.4167, 281.4568, 281.4971, 281.5374, 
    281.5774, 281.5461, 281.4719, 281.3975, 281.3232, 281.249, 281.1746, 
    281.1003, 281.0259, 280.9517, 280.8774, 280.803, 280.7288, 280.6545, 
    280.5801, 280.5251, 280.4854, 280.4456, 280.4058, 280.366, 280.3262, 
    280.2861, 280.2463, 280.2065, 280.1667, 280.127, 280.0872, 280.0474, 
    280.0076, 280.0234, 280.095, 280.1667, 280.2383, 280.3101, 280.3816, 
    280.4531, 280.5249, 280.5964, 280.6682, 280.7397, 280.8115, 280.8831, 
    280.9548, 280.9727, 280.9211, 280.8696, 280.8181, 280.7666, 280.7153, 
    280.6638, 280.6123, 280.5608, 280.5095, 280.458, 280.4065, 280.355, 
    280.3037, 280.2583, 280.2229, 280.1877, 280.1526, 280.1172, 280.082, 
    280.0469, 280.0117, 279.9763, 279.9412, 279.906, 279.8706, 279.8354, 
    279.8003, 279.7859, 279.8181, 279.8501, 279.8821, 279.9143, 279.9463, 
    279.9783, 280.0105, 280.0425, 280.0745, 280.1064, 280.1387, 280.1707, 
    280.2026, 280.2173, 280.1794, 280.1416, 280.1038, 280.0659, 280.0281, 
    279.9902, 279.9524, 279.9146, 279.8767, 279.8389, 279.801, 279.7632, 
    279.7253, 279.6821, 279.6165, 279.5505, 279.4846, 279.4187, 279.3528, 
    279.2869, 279.2212, 279.1553, 279.0894, 279.0234, 278.9575, 278.8916, 
    278.8259, 278.7639, 278.73, 278.6963, 278.6624, 278.6287, 278.5947, 
    278.5608, 278.5271, 278.4932, 278.4592, 278.4255, 278.3916, 278.3577, 
    278.324, 278.2927, 278.3003, 278.3079, 278.3157, 278.3232, 278.3311, 
    278.3386, 278.3462, 278.354, 278.3616, 278.3691, 278.377, 278.3845, 
    278.3921, 278.3999, 278.4053, 278.4109, 278.4163, 278.4216, 278.4272, 
    278.4326, 278.4382, 278.4436, 278.4492, 278.4546, 278.46, 278.4656, 
    278.4709, 278.4766, 278.4297, 278.3794, 278.3291, 278.2788, 278.2285, 
    278.1782, 278.1279, 278.0776, 278.0273, 277.9771, 277.9268,
  274.896, 274.9126, 274.9294, 274.946, 274.9629, 274.9795, 274.9963, 
    275.0171, 275.0649, 275.113, 275.1609, 275.209, 275.2568, 275.3049, 
    275.3528, 275.4009, 275.4487, 275.4968, 275.5447, 275.5928, 275.6406, 
    275.6924, 275.7986, 275.905, 276.0112, 276.1177, 276.2241, 276.3303, 
    276.4368, 276.543, 276.6494, 276.7556, 276.8621, 276.9685, 277.0747, 
    277.1812, 277.2637, 277.3462, 277.4287, 277.5112, 277.594, 277.6765, 
    277.759, 277.8416, 277.9241, 278.0066, 278.0891, 278.1719, 278.2544, 
    278.3369, 278.3198, 278.2959, 278.2722, 278.2485, 278.2246, 278.2009, 
    278.177, 278.1533, 278.1294, 278.1057, 278.082, 278.0581, 278.0344, 
    278.0105, 278.0427, 278.0828, 278.123, 278.1631, 278.2031, 278.2432, 
    278.2834, 278.3235, 278.3635, 278.4036, 278.4438, 278.4839, 278.5239, 
    278.5642, 278.6389, 278.7219, 278.8047, 278.8877, 278.9705, 279.0532, 
    279.1362, 279.219, 279.302, 279.3848, 279.4678, 279.5505, 279.6335, 
    279.7163, 279.804, 279.8931, 279.9822, 280.0713, 280.1606, 280.2498, 
    280.3389, 280.428, 280.5171, 280.6064, 280.6956, 280.7847, 280.8738, 
    280.9629, 281.0303, 281.0876, 281.145, 281.2024, 281.2598, 281.3171, 
    281.3745, 281.4319, 281.489, 281.5464, 281.6038, 281.6611, 281.7185, 
    281.7759, 281.7524, 281.6807, 281.6089, 281.5371, 281.4653, 281.3936, 
    281.3218, 281.25, 281.1782, 281.1064, 281.0347, 280.9629, 280.8911, 
    280.8193, 280.7581, 280.7051, 280.6519, 280.5986, 280.5457, 280.4924, 
    280.4395, 280.3862, 280.333, 280.28, 280.2268, 280.1736, 280.1206, 
    280.0674, 280.0784, 280.1533, 280.2285, 280.3035, 280.3784, 280.4536, 
    280.5286, 280.6035, 280.6787, 280.7537, 280.8286, 280.9036, 280.9788, 
    281.0537, 281.0759, 281.0298, 280.9839, 280.9377, 280.8918, 280.8459, 
    280.7998, 280.7539, 280.708, 280.6619, 280.616, 280.5701, 280.5239, 
    280.478, 280.4351, 280.397, 280.3589, 280.3208, 280.283, 280.2449, 
    280.2068, 280.1687, 280.1306, 280.0928, 280.0547, 280.0166, 279.9785, 
    279.9404, 279.9224, 279.948, 279.9736, 279.9993, 280.0249, 280.0505, 
    280.0764, 280.1021, 280.1277, 280.1533, 280.179, 280.2046, 280.2302, 
    280.2559, 280.2649, 280.2241, 280.1836, 280.1428, 280.1021, 280.0613, 
    280.0205, 279.9797, 279.9392, 279.8984, 279.8577, 279.8169, 279.7761, 
    279.7354, 279.6909, 279.6299, 279.5688, 279.5081, 279.447, 279.386, 
    279.325, 279.2639, 279.2029, 279.1418, 279.0811, 279.02, 278.959, 
    278.8979, 278.8396, 278.7988, 278.7583, 278.7178, 278.677, 278.6365, 
    278.5959, 278.5552, 278.5146, 278.4741, 278.4333, 278.3928, 278.3523, 
    278.3118, 278.2742, 278.2825, 278.291, 278.2993, 278.3079, 278.3162, 
    278.3247, 278.333, 278.3416, 278.3499, 278.3584, 278.3667, 278.3752, 
    278.3835, 278.3921, 278.4001, 278.4082, 278.4163, 278.4246, 278.4326, 
    278.4407, 278.4487, 278.4568, 278.4651, 278.4731, 278.4812, 278.4893, 
    278.4973, 278.5056, 278.4556, 278.4016, 278.3477, 278.2937, 278.2397, 
    278.1858, 278.1321, 278.0781, 278.0242, 277.9702, 277.9163,
  274.8938, 274.9155, 274.937, 274.9587, 274.9805, 275.002, 275.0237, 
    275.0476, 275.0869, 275.1262, 275.1655, 275.2048, 275.2441, 275.2834, 
    275.3228, 275.3621, 275.4014, 275.4407, 275.48, 275.5193, 275.5586, 
    275.6011, 275.6917, 275.7822, 275.8728, 275.9634, 276.054, 276.1445, 
    276.2351, 276.3257, 276.4163, 276.5068, 276.5974, 276.688, 276.7788, 
    276.8694, 276.9663, 277.0635, 277.1606, 277.2576, 277.3547, 277.4519, 
    277.5488, 277.646, 277.7429, 277.8401, 277.9373, 278.0342, 278.1313, 
    278.2285, 278.2314, 278.228, 278.2246, 278.2214, 278.218, 278.2146, 
    278.2112, 278.208, 278.2046, 278.2012, 278.198, 278.1946, 278.1912, 
    278.1877, 278.2214, 278.2605, 278.2993, 278.3381, 278.3772, 278.416, 
    278.4551, 278.4939, 278.533, 278.5718, 278.6106, 278.6497, 278.6885, 
    278.7275, 278.7942, 278.8672, 278.9402, 279.0134, 279.0864, 279.1594, 
    279.2327, 279.3057, 279.3787, 279.4517, 279.5249, 279.5979, 279.6709, 
    279.7441, 279.8259, 279.9106, 279.9956, 280.0803, 280.165, 280.25, 
    280.3347, 280.4194, 280.5044, 280.5891, 280.6738, 280.7585, 280.8435, 
    280.9282, 281.0059, 281.0803, 281.155, 281.2295, 281.304, 281.3784, 
    281.4529, 281.5273, 281.6018, 281.6763, 281.7507, 281.8252, 281.8997, 
    281.9744, 281.959, 281.8896, 281.8203, 281.7512, 281.6819, 281.6125, 
    281.5435, 281.4741, 281.4048, 281.3357, 281.2664, 281.1973, 281.1279, 
    281.0586, 280.991, 280.9246, 280.8582, 280.7917, 280.7253, 280.6589, 
    280.5925, 280.5261, 280.4595, 280.3931, 280.3267, 280.2603, 280.1938, 
    280.1274, 280.1335, 280.2119, 280.2903, 280.3687, 280.447, 280.5254, 
    280.6038, 280.6824, 280.7607, 280.8391, 280.9175, 280.9958, 281.0742, 
    281.1526, 281.179, 281.1387, 281.0981, 281.0576, 281.0171, 280.9766, 
    280.936, 280.8955, 280.855, 280.8145, 280.7739, 280.7334, 280.6929, 
    280.6526, 280.6118, 280.571, 280.53, 280.4893, 280.4485, 280.4077, 
    280.3667, 280.3259, 280.2852, 280.2441, 280.2034, 280.1626, 280.1216, 
    280.0808, 280.0588, 280.0781, 280.0972, 280.1165, 280.1357, 280.155, 
    280.1743, 280.1936, 280.2129, 280.2319, 280.2512, 280.2705, 280.2898, 
    280.3091, 280.3125, 280.269, 280.2253, 280.1816, 280.1382, 280.0945, 
    280.0508, 280.0073, 279.9636, 279.9202, 279.8765, 279.8328, 279.7893, 
    279.7456, 279.6997, 279.6436, 279.5874, 279.5312, 279.4751, 279.4189, 
    279.363, 279.3069, 279.2507, 279.1946, 279.1384, 279.0823, 279.0261, 
    278.9702, 278.915, 278.8677, 278.8203, 278.7729, 278.7256, 278.6782, 
    278.6309, 278.5835, 278.5361, 278.4888, 278.4414, 278.394, 278.3467, 
    278.2993, 278.2556, 278.2646, 278.2739, 278.2832, 278.2922, 278.3015, 
    278.3108, 278.3198, 278.3291, 278.3384, 278.3474, 278.3567, 278.366, 
    278.375, 278.3843, 278.395, 278.4058, 278.4165, 278.4272, 278.438, 
    278.4487, 278.4595, 278.4702, 278.481, 278.4917, 278.5024, 278.5132, 
    278.5239, 278.5344, 278.4812, 278.4238, 278.3662, 278.3086, 278.2512, 
    278.1936, 278.136, 278.0786, 278.021, 277.9634, 277.906,
  274.9866, 275.0098, 275.033, 275.0559, 275.0791, 275.1023, 275.1255, 
    275.1514, 275.196, 275.241, 275.2856, 275.3306, 275.3752, 275.4202, 
    275.4648, 275.5098, 275.5544, 275.5994, 275.644, 275.689, 275.7336, 
    275.7805, 275.8584, 275.9365, 276.0144, 276.0925, 276.1704, 276.2485, 
    276.3264, 276.4045, 276.4824, 276.5605, 276.6384, 276.7163, 276.7944, 
    276.8723, 276.9556, 277.0386, 277.1216, 277.2046, 277.2876, 277.3706, 
    277.4539, 277.5369, 277.6199, 277.7029, 277.7859, 277.8691, 277.9521, 
    278.0352, 278.0554, 278.0713, 278.0874, 278.1035, 278.1194, 278.1355, 
    278.1514, 278.1675, 278.1836, 278.1995, 278.2156, 278.2314, 278.2476, 
    278.2637, 278.3081, 278.3564, 278.405, 278.4536, 278.502, 278.5505, 
    278.5991, 278.6475, 278.696, 278.7446, 278.793, 278.8416, 278.8899, 
    278.9385, 279.0007, 279.0659, 279.1311, 279.1963, 279.2617, 279.3269, 
    279.3921, 279.4573, 279.5227, 279.5879, 279.6531, 279.7185, 279.7837, 
    279.8489, 279.9253, 280.0054, 280.0852, 280.1653, 280.2454, 280.3254, 
    280.4055, 280.4856, 280.5654, 280.6455, 280.7256, 280.8057, 280.8857, 
    280.9658, 281.0447, 281.1233, 281.2019, 281.2805, 281.3591, 281.4377, 
    281.5164, 281.595, 281.6733, 281.752, 281.8306, 281.9092, 281.9878, 
    282.0664, 282.0557, 281.9907, 281.9248, 281.8579, 281.7903, 281.7214, 
    281.6516, 281.5808, 281.509, 281.4363, 281.3621, 281.2871, 281.2109, 
    281.1333, 281.0627, 280.9985, 280.9353, 280.873, 280.8118, 280.7515, 
    280.6919, 280.6333, 280.5754, 280.5186, 280.4624, 280.407, 280.3523, 
    280.2986, 280.3069, 280.3772, 280.4475, 280.5178, 280.5879, 280.6582, 
    280.7285, 280.7988, 280.8691, 280.9392, 281.0095, 281.0798, 281.1501, 
    281.2202, 281.2432, 281.2051, 281.167, 281.1292, 281.0911, 281.053, 
    281.0149, 280.9768, 280.9387, 280.9009, 280.8628, 280.8247, 280.7866, 
    280.7485, 280.71, 280.6699, 280.6301, 280.5901, 280.5503, 280.5105, 
    280.4705, 280.4307, 280.3909, 280.3508, 280.311, 280.2712, 280.2312, 
    280.1914, 280.1682, 280.1821, 280.1958, 280.2095, 280.2234, 280.2371, 
    280.2507, 280.2644, 280.2783, 280.292, 280.3057, 280.3196, 280.3333, 
    280.3469, 280.3464, 280.303, 280.2595, 280.2161, 280.1726, 280.1292, 
    280.0857, 280.0422, 279.9988, 279.9553, 279.9119, 279.8684, 279.825, 
    279.7815, 279.7361, 279.6819, 279.6274, 279.5732, 279.5188, 279.4646, 
    279.4104, 279.356, 279.3018, 279.2473, 279.1931, 279.1387, 279.0845, 
    279.0303, 278.9761, 278.9236, 278.8713, 278.8188, 278.7664, 278.7139, 
    278.6614, 278.6089, 278.5566, 278.5042, 278.4517, 278.3992, 278.3467, 
    278.2944, 278.2456, 278.2532, 278.2607, 278.2681, 278.2756, 278.2832, 
    278.2908, 278.2981, 278.3057, 278.3132, 278.3208, 278.3281, 278.3357, 
    278.3433, 278.3508, 278.3643, 278.3779, 278.3914, 278.4048, 278.4185, 
    278.4319, 278.4453, 278.459, 278.4724, 278.4858, 278.4995, 278.5129, 
    278.5264, 278.54, 278.4976, 278.4514, 278.4055, 278.3594, 278.3132, 
    278.2671, 278.2212, 278.175, 278.1289, 278.0828, 278.0366,
  275.0952, 275.1194, 275.1433, 275.1675, 275.1917, 275.2156, 275.2397, 
    275.2673, 275.3201, 275.3728, 275.4253, 275.478, 275.5308, 275.5833, 
    275.636, 275.6887, 275.7412, 275.7939, 275.8467, 275.8992, 275.9519, 
    276.0054, 276.0713, 276.1372, 276.2031, 276.269, 276.335, 276.4009, 
    276.4668, 276.5327, 276.5986, 276.6646, 276.7305, 276.7964, 276.8623, 
    276.9282, 276.9924, 277.0566, 277.1211, 277.1853, 277.2495, 277.3137, 
    277.3779, 277.4421, 277.5063, 277.5706, 277.635, 277.6992, 277.7634, 
    277.8276, 277.8647, 277.8999, 277.9351, 277.9702, 278.0054, 278.0408, 
    278.0759, 278.1111, 278.1462, 278.1814, 278.2168, 278.252, 278.2871, 
    278.3223, 278.3792, 278.439, 278.4988, 278.5588, 278.6187, 278.6785, 
    278.7385, 278.7983, 278.8582, 278.918, 278.978, 279.0378, 279.0977, 
    279.1575, 279.2158, 279.2734, 279.3313, 279.3889, 279.4468, 279.5046, 
    279.5623, 279.6201, 279.6777, 279.7356, 279.7935, 279.8511, 279.9089, 
    279.9666, 280.0376, 280.1128, 280.188, 280.2632, 280.3384, 280.4136, 
    280.4888, 280.564, 280.6392, 280.7144, 280.7896, 280.865, 280.9402, 
    281.0154, 281.0942, 281.1746, 281.2551, 281.3357, 281.4163, 281.4966, 
    281.5771, 281.6577, 281.7383, 281.8186, 281.8992, 281.9797, 282.0603, 
    282.1406, 282.1348, 282.0757, 282.0149, 281.9519, 281.8872, 281.8201, 
    281.7507, 281.6792, 281.6052, 281.5286, 281.449, 281.3667, 281.2815, 
    281.1929, 281.1187, 281.0596, 281.0027, 280.9475, 280.8945, 280.8433, 
    280.7939, 280.7461, 280.6997, 280.655, 280.6118, 280.5698, 280.5291, 
    280.4895, 280.5002, 280.5605, 280.6206, 280.6809, 280.741, 280.8013, 
    280.8613, 280.9216, 280.9817, 281.042, 281.1021, 281.1624, 281.2224, 
    281.2827, 281.3008, 281.2646, 281.2285, 281.1924, 281.1562, 281.1204, 
    281.0842, 281.0481, 281.012, 280.9758, 280.9399, 280.9038, 280.8677, 
    280.8315, 280.7947, 280.7563, 280.718, 280.6797, 280.6416, 280.6033, 
    280.5649, 280.5266, 280.4885, 280.4502, 280.4119, 280.3735, 280.3352, 
    280.2971, 280.2734, 280.2817, 280.29, 280.2986, 280.3069, 280.3152, 
    280.3237, 280.332, 280.3406, 280.3489, 280.3572, 280.3657, 280.374, 
    280.3823, 280.3779, 280.3352, 280.2925, 280.2498, 280.2068, 280.1641, 
    280.1213, 280.0786, 280.0359, 279.9929, 279.9502, 279.9075, 279.8647, 
    279.8218, 279.7771, 279.7241, 279.6711, 279.6182, 279.5652, 279.5122, 
    279.4592, 279.4062, 279.3533, 279.3003, 279.2473, 279.1943, 279.1411, 
    279.0881, 279.0347, 278.9775, 278.9202, 278.863, 278.8057, 278.7485, 
    278.6912, 278.634, 278.5767, 278.5195, 278.4622, 278.405, 278.3477, 
    278.2905, 278.2371, 278.2427, 278.248, 278.2534, 278.2588, 278.2642, 
    278.2695, 278.2751, 278.2805, 278.2859, 278.2913, 278.2966, 278.3022, 
    278.3076, 278.313, 278.3293, 278.3457, 278.3621, 278.3782, 278.3945, 
    278.4109, 278.4272, 278.4436, 278.46, 278.4761, 278.4924, 278.5088, 
    278.5251, 278.5415, 278.5125, 278.4802, 278.4482, 278.416, 278.3838, 
    278.3518, 278.3196, 278.2876, 278.2554, 278.2234, 278.1912,
  275.2039, 275.2288, 275.2539, 275.2788, 275.304, 275.3289, 275.354, 
    275.3833, 275.4438, 275.5044, 275.5649, 275.6255, 275.686, 275.7466, 
    275.8071, 275.8677, 275.928, 275.9885, 276.0491, 276.1096, 276.1702, 
    276.2302, 276.2842, 276.3379, 276.3918, 276.4456, 276.4995, 276.5535, 
    276.6072, 276.6611, 276.7148, 276.7688, 276.8225, 276.8765, 276.9302, 
    276.9841, 277.0295, 277.075, 277.1204, 277.1658, 277.2112, 277.2566, 
    277.302, 277.3477, 277.3931, 277.4385, 277.4839, 277.5293, 277.5747, 
    277.6201, 277.6738, 277.7283, 277.7827, 277.8372, 277.8916, 277.9458, 
    278.0002, 278.0547, 278.1091, 278.1636, 278.2178, 278.2722, 278.3267, 
    278.3811, 278.4502, 278.5215, 278.5928, 278.6641, 278.7354, 278.8066, 
    278.8777, 278.949, 279.0203, 279.0916, 279.1628, 279.2341, 279.3054, 
    279.3767, 279.4309, 279.4812, 279.5315, 279.5818, 279.6318, 279.6821, 
    279.7324, 279.7827, 279.833, 279.8833, 279.9336, 279.9839, 280.0342, 
    280.0845, 280.1497, 280.2202, 280.2905, 280.3608, 280.4314, 280.5017, 
    280.572, 280.6426, 280.7129, 280.7832, 280.8538, 280.9241, 280.9944, 
    281.0649, 281.1436, 281.2261, 281.3083, 281.3909, 281.4731, 281.5557, 
    281.6379, 281.7205, 281.803, 281.8853, 281.9678, 282.05, 282.1326, 
    282.2151, 282.2148, 282.1631, 282.1089, 282.052, 281.9922, 281.9292, 
    281.8625, 281.7922, 281.718, 281.6394, 281.5557, 281.467, 281.3723, 
    281.2712, 281.1926, 281.1379, 281.0869, 281.0388, 280.9937, 280.9512, 
    280.9109, 280.8728, 280.8369, 280.8027, 280.7703, 280.7395, 280.7102, 
    280.6821, 280.6936, 280.7439, 280.7939, 280.844, 280.894, 280.9443, 
    280.9944, 281.0444, 281.0945, 281.1445, 281.1948, 281.2449, 281.2949, 
    281.345, 281.3582, 281.3242, 281.29, 281.2559, 281.2217, 281.1875, 
    281.1536, 281.1194, 281.0852, 281.051, 281.0168, 280.9829, 280.9487, 
    280.9146, 280.8794, 280.8428, 280.8062, 280.7693, 280.7327, 280.696, 
    280.6594, 280.6228, 280.5859, 280.5493, 280.5127, 280.4761, 280.4392, 
    280.4026, 280.3784, 280.3813, 280.3845, 280.3875, 280.3906, 280.3936, 
    280.3965, 280.3997, 280.4026, 280.4058, 280.4087, 280.4119, 280.4148, 
    280.4177, 280.4097, 280.3674, 280.3254, 280.2832, 280.2412, 280.199, 
    280.157, 280.1147, 280.0728, 280.0305, 279.9885, 279.9463, 279.9043, 
    279.8621, 279.8184, 279.7666, 279.7148, 279.6631, 279.6116, 279.5598, 
    279.5081, 279.4565, 279.4048, 279.353, 279.3013, 279.2498, 279.198, 
    279.1462, 279.0933, 279.0312, 278.9692, 278.9072, 278.8452, 278.783, 
    278.7209, 278.6589, 278.5969, 278.5349, 278.4729, 278.4106, 278.3486, 
    278.2866, 278.2288, 278.2319, 278.2354, 278.2388, 278.2419, 278.2454, 
    278.2485, 278.252, 278.2554, 278.2585, 278.262, 278.2651, 278.2686, 
    278.272, 278.2751, 278.2944, 278.3135, 278.3325, 278.3518, 278.3708, 
    278.3899, 278.4092, 278.4282, 278.4473, 278.4666, 278.4856, 278.5046, 
    278.5239, 278.543, 278.5271, 278.509, 278.491, 278.4727, 278.4546, 
    278.4365, 278.4182, 278.4001, 278.3821, 278.3638, 278.3457,
  275.3125, 275.3384, 275.3645, 275.3904, 275.4163, 275.4421, 275.4683, 
    275.4995, 275.5679, 275.6362, 275.7046, 275.7729, 275.8413, 275.9097, 
    275.978, 276.0466, 276.115, 276.1833, 276.2517, 276.3201, 276.3884, 
    276.4551, 276.4968, 276.5388, 276.5806, 276.6223, 276.6641, 276.7058, 
    276.7476, 276.7893, 276.8311, 276.8728, 276.9146, 276.9563, 276.9983, 
    277.04, 277.0667, 277.0933, 277.1199, 277.1465, 277.1731, 277.1997, 
    277.2263, 277.2529, 277.2795, 277.3062, 277.3328, 277.3594, 277.386, 
    277.4126, 277.4832, 277.5569, 277.6304, 277.7041, 277.7776, 277.8511, 
    277.9248, 277.9983, 278.0718, 278.1455, 278.219, 278.2927, 278.3662, 
    278.4397, 278.5212, 278.604, 278.6865, 278.7693, 278.8518, 278.9346, 
    279.0171, 279.0999, 279.1824, 279.2651, 279.3477, 279.4304, 279.5129, 
    279.5957, 279.646, 279.6887, 279.7314, 279.7744, 279.8171, 279.8599, 
    279.9026, 279.9456, 279.9883, 280.031, 280.0737, 280.1167, 280.1594, 
    280.2021, 280.262, 280.3276, 280.3931, 280.4587, 280.5244, 280.5898, 
    280.6555, 280.7209, 280.7866, 280.8523, 280.9177, 280.9834, 281.0488, 
    281.1145, 281.1929, 281.2773, 281.3616, 281.446, 281.5303, 281.6145, 
    281.699, 281.7832, 281.8677, 281.9519, 282.0364, 282.1206, 282.2051, 
    282.2893, 282.2957, 282.2529, 282.2075, 282.1587, 282.1064, 282.05, 
    281.9895, 281.9238, 281.8525, 281.7749, 281.6899, 281.5967, 281.4939, 
    281.3799, 281.2944, 281.2424, 281.1956, 281.1531, 281.1143, 281.0789, 
    281.0464, 281.0164, 280.9888, 280.9629, 280.939, 280.9167, 280.896, 
    280.8765, 280.887, 280.927, 280.967, 281.0071, 281.0471, 281.0872, 
    281.1272, 281.1672, 281.2073, 281.2473, 281.2874, 281.3274, 281.3674, 
    281.4075, 281.4158, 281.3835, 281.3516, 281.3193, 281.2871, 281.2549, 
    281.2227, 281.1907, 281.1584, 281.1262, 281.094, 281.0618, 281.0298, 
    280.9976, 280.9644, 280.9292, 280.894, 280.8591, 280.824, 280.7888, 
    280.7537, 280.7188, 280.6836, 280.6484, 280.6135, 280.5784, 280.5432, 
    280.5083, 280.4834, 280.481, 280.4788, 280.4766, 280.4741, 280.4719, 
    280.4695, 280.4673, 280.4648, 280.4626, 280.4602, 280.458, 280.4556, 
    280.4534, 280.4412, 280.3997, 280.3584, 280.3169, 280.2754, 280.2339, 
    280.1926, 280.1511, 280.1096, 280.0681, 280.0269, 279.9854, 279.9438, 
    279.9026, 279.8594, 279.8091, 279.7585, 279.7083, 279.6577, 279.6074, 
    279.5571, 279.5066, 279.4563, 279.4058, 279.3555, 279.3052, 279.2546, 
    279.2043, 279.1519, 279.085, 279.0181, 278.9514, 278.8845, 278.8176, 
    278.7507, 278.6838, 278.6172, 278.5503, 278.4834, 278.4165, 278.3496, 
    278.2827, 278.2202, 278.2214, 278.2227, 278.2239, 278.2251, 278.2263, 
    278.2275, 278.2288, 278.23, 278.2312, 278.2324, 278.2336, 278.2349, 
    278.2361, 278.2373, 278.2593, 278.2812, 278.3032, 278.3252, 278.3472, 
    278.3689, 278.3909, 278.4128, 278.4348, 278.4568, 278.4788, 278.5005, 
    278.5225, 278.5444, 278.542, 278.5378, 278.5334, 278.5293, 278.5251, 
    278.521, 278.5168, 278.5127, 278.5085, 278.5044, 278.5002,
  275.4211, 275.448, 275.4749, 275.5017, 275.5286, 275.5557, 275.5825, 
    275.6155, 275.6917, 275.7681, 275.8442, 275.9204, 275.9968, 276.073, 
    276.1492, 276.2256, 276.3018, 276.3779, 276.4541, 276.5305, 276.6067, 
    276.6802, 276.7097, 276.7395, 276.769, 276.7988, 276.8286, 276.8582, 
    276.8879, 276.9177, 276.9473, 276.9771, 277.0068, 277.0364, 277.0662, 
    277.0957, 277.1035, 277.1113, 277.1191, 277.127, 277.1348, 277.1426, 
    277.1504, 277.1582, 277.166, 277.1738, 277.1816, 277.1895, 277.1973, 
    277.2051, 277.2925, 277.3853, 277.478, 277.5708, 277.6636, 277.7563, 
    277.8491, 277.9419, 278.0347, 278.1274, 278.2202, 278.313, 278.4058, 
    278.4985, 278.5923, 278.6865, 278.7805, 278.8745, 278.9685, 279.0625, 
    279.1565, 279.2505, 279.3447, 279.4387, 279.5327, 279.6267, 279.7207, 
    279.8147, 279.8611, 279.8965, 279.9316, 279.967, 280.0022, 280.0376, 
    280.0728, 280.1082, 280.1433, 280.1787, 280.2141, 280.2493, 280.2847, 
    280.3198, 280.3743, 280.4351, 280.4958, 280.5566, 280.6172, 280.678, 
    280.7388, 280.7996, 280.8604, 280.9211, 280.9817, 281.0425, 281.1033, 
    281.1641, 281.2424, 281.3286, 281.4148, 281.501, 281.5874, 281.6736, 
    281.7598, 281.8462, 281.9324, 282.0186, 282.105, 282.1912, 282.2773, 
    282.3635, 282.3772, 282.3452, 282.3105, 282.2727, 282.231, 282.1853, 
    282.1348, 282.0784, 282.0154, 281.9443, 281.8638, 281.7715, 281.6648, 
    281.54, 281.4434, 281.3884, 281.3413, 281.3005, 281.2646, 281.2332, 
    281.2053, 281.1802, 281.1577, 281.1372, 281.1189, 281.1018, 281.0864, 
    281.0723, 281.0806, 281.1104, 281.1404, 281.1704, 281.2002, 281.2302, 
    281.26, 281.29, 281.3201, 281.3499, 281.3799, 281.4099, 281.4397, 
    281.4697, 281.4734, 281.4431, 281.4128, 281.3828, 281.3525, 281.3223, 
    281.292, 281.2617, 281.2317, 281.2014, 281.1711, 281.1409, 281.1106, 
    281.0806, 281.0491, 281.0156, 280.9822, 280.9487, 280.915, 280.8816, 
    280.8481, 280.8147, 280.7812, 280.7478, 280.7144, 280.6809, 280.6472, 
    280.6138, 280.5884, 280.5808, 280.573, 280.5654, 280.5576, 280.55, 
    280.5425, 280.5347, 280.5271, 280.5193, 280.5117, 280.5039, 280.4963, 
    280.4888, 280.4727, 280.4319, 280.3911, 280.3503, 280.3096, 280.2688, 
    280.228, 280.1873, 280.1465, 280.106, 280.0652, 280.0244, 279.9836, 
    279.9429, 279.9004, 279.8513, 279.8022, 279.7532, 279.7041, 279.655, 
    279.606, 279.5569, 279.5078, 279.4587, 279.4097, 279.3606, 279.3115, 
    279.2625, 279.2104, 279.1389, 279.0671, 278.9956, 278.9238, 278.8523, 
    278.7805, 278.709, 278.6372, 278.5657, 278.4939, 278.4224, 278.3506, 
    278.2791, 278.2117, 278.2109, 278.21, 278.2092, 278.2083, 278.2075, 
    278.2065, 278.2056, 278.2048, 278.2039, 278.2031, 278.2021, 278.2014, 
    278.2004, 278.1997, 278.2244, 278.249, 278.2739, 278.2986, 278.3232, 
    278.3481, 278.3728, 278.3975, 278.4224, 278.447, 278.4717, 278.4966, 
    278.5212, 278.5459, 278.5566, 278.5664, 278.5762, 278.5862, 278.5959, 
    278.6057, 278.6155, 278.6252, 278.635, 278.6448, 278.6545,
  275.5298, 275.5576, 275.5854, 275.6133, 275.6411, 275.6689, 275.6965, 
    275.7314, 275.8157, 275.8997, 275.9839, 276.0679, 276.1521, 276.2361, 
    276.3203, 276.4043, 276.4885, 276.5728, 276.6567, 276.741, 276.825, 
    276.905, 276.9226, 276.9402, 276.9578, 276.9753, 276.9932, 277.0107, 
    277.0283, 277.0459, 277.0635, 277.0813, 277.0989, 277.1165, 277.134, 
    277.1516, 277.1406, 277.1296, 277.1187, 277.1077, 277.0967, 277.0857, 
    277.0747, 277.0637, 277.0525, 277.0415, 277.0305, 277.0195, 277.0085, 
    276.9976, 277.1018, 277.2139, 277.3257, 277.4377, 277.5496, 277.6616, 
    277.7737, 277.8855, 277.9976, 278.1094, 278.2214, 278.3333, 278.4453, 
    278.5574, 278.6636, 278.7688, 278.8743, 278.9797, 279.0852, 279.1904, 
    279.2959, 279.4014, 279.5068, 279.6123, 279.7175, 279.823, 279.9285, 
    280.0339, 280.0762, 280.104, 280.1318, 280.1597, 280.1875, 280.2153, 
    280.2429, 280.2708, 280.2986, 280.3264, 280.3542, 280.3821, 280.4099, 
    280.4377, 280.4866, 280.5425, 280.5984, 280.6543, 280.7102, 280.7661, 
    280.822, 280.8782, 280.9341, 280.99, 281.0459, 281.1018, 281.1577, 
    281.2136, 281.2917, 281.3799, 281.468, 281.5562, 281.6443, 281.7327, 
    281.8208, 281.9089, 281.9971, 282.0852, 282.1733, 282.2615, 282.3499, 
    282.438, 282.4597, 282.4402, 282.4187, 282.3948, 282.3677, 282.3372, 
    282.3025, 282.3755, 282.3713, 282.3677, 282.3647, 282.3621, 282.3596, 
    282.3577, 282.3464, 281.6069, 281.5466, 281.4976, 281.457, 281.4231, 
    281.394, 281.3689, 281.3472, 281.3279, 281.3108, 281.2957, 281.282, 
    281.2695, 281.2739, 281.2937, 281.3135, 281.3335, 281.3533, 281.373, 
    281.3931, 281.4128, 281.4329, 281.4526, 281.4724, 281.4924, 281.5122, 
    281.532, 281.531, 281.5027, 281.4744, 281.446, 281.4177, 281.3896, 
    281.3613, 281.333, 281.3047, 281.2766, 281.2483, 281.22, 281.1917, 
    281.1636, 281.1338, 281.1021, 281.0701, 281.0383, 281.0063, 280.9744, 
    280.9426, 280.9106, 280.8789, 280.8469, 280.8152, 280.7832, 280.7512, 
    280.7195, 280.6934, 280.6804, 280.6675, 280.6543, 280.6414, 280.6284, 
    280.6152, 280.6023, 280.5891, 280.5762, 280.5632, 280.55, 280.5371, 
    280.5242, 280.5044, 280.4641, 280.4241, 280.384, 280.344, 280.3037, 
    280.2637, 280.2236, 280.1836, 280.1436, 280.1033, 280.0632, 280.0232, 
    279.9832, 279.9417, 279.8938, 279.8459, 279.7981, 279.7505, 279.7026, 
    279.6548, 279.6072, 279.5593, 279.5115, 279.4639, 279.416, 279.3682, 
    279.3203, 279.269, 279.1926, 279.1162, 279.0398, 278.9631, 278.8867, 
    278.8103, 278.7339, 278.6575, 278.5811, 278.5044, 278.428, 278.3516, 
    278.2751, 278.2034, 278.2004, 278.1973, 278.1943, 278.1914, 278.1885, 
    278.1855, 278.1826, 278.1797, 278.1765, 278.1736, 278.1707, 278.1677, 
    278.1648, 278.1619, 278.1895, 278.2168, 278.2444, 278.272, 278.2996, 
    278.3271, 278.3547, 278.3821, 278.4097, 278.4373, 278.4648, 278.4924, 
    278.5198, 278.5474, 278.5715, 278.5952, 278.6189, 278.6428, 278.6665, 
    278.6902, 278.7141, 278.7378, 278.7615, 278.7854, 278.8091,
  275.6384, 275.6672, 275.696, 275.7246, 275.7534, 275.7822, 275.8108, 
    275.8474, 275.9395, 276.0315, 276.1235, 276.2153, 276.3074, 276.3994, 
    276.4915, 276.5833, 276.6753, 276.7673, 276.8594, 276.9512, 277.0432, 
    277.1299, 277.1355, 277.1409, 277.1465, 277.1521, 277.1575, 277.1631, 
    277.1687, 277.1743, 277.1797, 277.1853, 277.1909, 277.1965, 277.2019, 
    277.2075, 277.1777, 277.1479, 277.1182, 277.0881, 277.0583, 277.0286, 
    276.9988, 276.969, 276.9392, 276.9094, 276.8794, 276.8496, 276.8198, 
    276.79, 276.9111, 277.0422, 277.1733, 277.3044, 277.4358, 277.5669, 
    277.698, 277.8291, 277.9602, 278.0913, 278.2227, 278.3538, 278.4849, 
    278.616, 278.7346, 278.8513, 278.9683, 279.085, 279.2017, 279.3186, 
    279.4353, 279.5522, 279.6689, 279.7856, 279.9026, 280.0193, 280.136, 
    280.2529, 280.2913, 280.3115, 280.332, 280.3523, 280.3726, 280.3928, 
    280.4131, 280.4336, 280.4539, 280.4741, 280.4944, 280.5149, 280.5352, 
    280.5554, 280.5989, 280.6499, 280.7009, 280.7522, 280.8032, 280.8542, 
    280.9055, 280.9565, 281.0076, 281.0588, 281.1099, 281.1609, 281.2122, 
    281.2632, 281.3411, 281.4312, 281.5212, 281.6113, 281.7014, 281.7915, 
    281.8816, 281.9717, 282.0618, 282.1519, 282.2419, 282.332, 282.4221, 
    282.5122, 282.5432, 282.5381, 282.5322, 282.5256, 282.5181, 282.5093, 
    282.499, 282.4231, 282.4182, 282.4143, 282.4106, 282.4077, 282.405, 
    282.4028, 282.3938, 281.9697, 281.8574, 281.7751, 281.7122, 281.6624, 
    281.6221, 281.5886, 281.5608, 281.5369, 281.5164, 281.4983, 281.4827, 
    281.4688, 281.4673, 281.4771, 281.4868, 281.4966, 281.5063, 281.5161, 
    281.5259, 281.5356, 281.5454, 281.5554, 281.5652, 281.575, 281.5847, 
    281.5945, 281.5884, 281.5623, 281.5359, 281.5095, 281.4832, 281.4568, 
    281.4307, 281.4043, 281.3779, 281.3516, 281.3254, 281.2991, 281.2727, 
    281.2463, 281.2188, 281.1885, 281.1582, 281.1279, 281.0977, 281.0674, 
    281.0371, 281.0066, 280.9763, 280.946, 280.9158, 280.8855, 280.8552, 
    280.825, 280.7986, 280.78, 280.7617, 280.7434, 280.7249, 280.7065, 
    280.6882, 280.6699, 280.6514, 280.6331, 280.6147, 280.5962, 280.5779, 
    280.5596, 280.5359, 280.4963, 280.457, 280.4175, 280.3782, 280.3389, 
    280.2993, 280.26, 280.2205, 280.1812, 280.1416, 280.1023, 280.0627, 
    280.0234, 279.9827, 279.9363, 279.8896, 279.8433, 279.7966, 279.7502, 
    279.7039, 279.6572, 279.6108, 279.5645, 279.5178, 279.4714, 279.425, 
    279.3784, 279.3276, 279.2463, 279.165, 279.084, 279.0027, 278.9214, 
    278.8401, 278.7588, 278.6775, 278.5964, 278.5151, 278.4338, 278.3525, 
    278.2712, 278.1948, 278.1897, 278.1848, 278.1797, 278.1746, 278.1694, 
    278.1646, 278.1594, 278.1543, 278.1494, 278.1443, 278.1392, 278.134, 
    278.1292, 278.124, 278.1543, 278.1848, 278.2151, 278.2454, 278.2759, 
    278.3062, 278.3364, 278.3669, 278.3972, 278.4275, 278.4578, 278.4883, 
    278.5186, 278.5488, 278.5862, 278.624, 278.6616, 278.6995, 278.7371, 
    278.7749, 278.8127, 278.8503, 278.8882, 278.9258, 278.9636,
  275.8152, 275.8481, 275.8811, 275.9141, 275.947, 275.9802, 276.0132, 
    276.0537, 276.1484, 276.2432, 276.3379, 276.4326, 276.5273, 276.6221, 
    276.7168, 276.8115, 276.9062, 277.001, 277.0955, 277.1902, 277.2849, 
    277.3752, 277.3982, 277.4214, 277.4443, 277.4675, 277.4905, 277.5137, 
    277.5366, 277.5596, 277.5828, 277.6057, 277.6289, 277.6519, 277.675, 
    277.698, 277.6367, 277.5752, 277.5137, 277.4524, 277.3909, 277.3296, 
    277.2681, 277.2068, 277.1453, 277.084, 277.0225, 276.9612, 276.8997, 
    276.8384, 276.95, 277.0732, 277.1968, 277.3201, 277.4434, 277.5667, 
    277.6899, 277.8132, 277.9365, 278.0598, 278.1831, 278.3066, 278.4299, 
    278.5532, 278.6768, 278.8005, 278.9243, 279.0479, 279.1716, 279.2952, 
    279.4189, 279.5427, 279.6663, 279.79, 279.9138, 280.0374, 280.1611, 
    280.2849, 280.3271, 280.3511, 280.3748, 280.3984, 280.4221, 280.4458, 
    280.4695, 280.4932, 280.5168, 280.5405, 280.5645, 280.5881, 280.6118, 
    280.6355, 280.677, 280.7241, 280.7715, 280.8188, 280.8662, 280.9136, 
    280.9609, 281.0083, 281.0557, 281.1028, 281.1501, 281.1975, 281.2449, 
    281.2922, 281.3628, 281.4441, 281.5251, 281.6064, 281.6875, 281.7688, 
    281.8499, 281.9312, 282.0122, 282.0935, 282.1748, 282.2559, 282.3372, 
    282.4182, 282.4441, 282.436, 282.427, 282.417, 282.4055, 282.3926, 
    282.3777, 282.3984, 282.3962, 282.3945, 282.3928, 282.3916, 282.3904, 
    282.3894, 282.3804, 281.9138, 281.8279, 281.7603, 281.7056, 281.6604, 
    281.6226, 281.5903, 281.5625, 281.5383, 281.5171, 281.4983, 281.4817, 
    281.4666, 281.4619, 281.4663, 281.4709, 281.4753, 281.48, 281.4844, 
    281.489, 281.4934, 281.4978, 281.5024, 281.5068, 281.5115, 281.5159, 
    281.5205, 281.5146, 281.4956, 281.4766, 281.4575, 281.4385, 281.4194, 
    281.4006, 281.3816, 281.3625, 281.3435, 281.3245, 281.3054, 281.2864, 
    281.2673, 281.2466, 281.2227, 281.1987, 281.1748, 281.1509, 281.127, 
    281.1033, 281.0793, 281.0554, 281.0315, 281.0076, 280.9836, 280.9597, 
    280.9358, 280.9111, 280.8845, 280.8577, 280.8311, 280.8042, 280.7776, 
    280.7507, 280.7241, 280.6973, 280.6707, 280.644, 280.6172, 280.5906, 
    280.5637, 280.5342, 280.4956, 280.4568, 280.4182, 280.3796, 280.3411, 
    280.3025, 280.2639, 280.2253, 280.1868, 280.1482, 280.1094, 280.0708, 
    280.0322, 279.9924, 279.9478, 279.9031, 279.8584, 279.8137, 279.769, 
    279.7244, 279.6797, 279.635, 279.5903, 279.5457, 279.501, 279.4563, 
    279.4116, 279.3628, 279.2834, 279.2041, 279.1248, 279.0454, 278.9661, 
    278.8867, 278.8074, 278.728, 278.6487, 278.5693, 278.49, 278.4106, 
    278.3313, 278.2563, 278.2478, 278.239, 278.2302, 278.2214, 278.2129, 
    278.2041, 278.1953, 278.1868, 278.178, 278.1692, 278.1604, 278.1519, 
    278.1431, 278.1343, 278.1631, 278.1917, 278.2205, 278.2493, 278.2778, 
    278.3066, 278.3354, 278.364, 278.3928, 278.4216, 278.4502, 278.479, 
    278.5078, 278.5364, 278.5686, 278.6011, 278.6335, 278.666, 278.6987, 
    278.7312, 278.7637, 278.7961, 278.8286, 278.8611, 278.8936,
  276.0061, 276.0439, 276.0818, 276.1199, 276.1577, 276.1956, 276.2336, 
    276.2788, 276.3752, 276.4714, 276.5679, 276.6643, 276.7607, 276.8569, 
    276.9534, 277.0498, 277.146, 277.2424, 277.3389, 277.4353, 277.5315, 
    277.6248, 277.6716, 277.7183, 277.7649, 277.8118, 277.8584, 277.905, 
    277.9519, 277.9985, 278.0452, 278.092, 278.1387, 278.1853, 278.2322, 
    278.2788, 278.1831, 278.0874, 277.9919, 277.8962, 277.8005, 277.7048, 
    277.6091, 277.5137, 277.418, 277.3223, 277.2266, 277.1309, 277.0352, 
    276.9397, 277.0366, 277.1465, 277.2563, 277.3662, 277.4761, 277.5859, 
    277.696, 277.8059, 277.9158, 278.0256, 278.1355, 278.2454, 278.3552, 
    278.4651, 278.5923, 278.7219, 278.8516, 278.9812, 279.1108, 279.2405, 
    279.3704, 279.5, 279.6296, 279.7593, 279.8889, 280.0186, 280.1482, 
    280.2778, 280.3259, 280.3555, 280.3848, 280.4141, 280.4434, 280.4729, 
    280.5022, 280.5315, 280.5608, 280.5903, 280.6196, 280.6489, 280.6782, 
    280.7078, 280.7478, 280.7917, 280.8354, 280.8792, 280.9229, 280.9668, 
    281.0105, 281.0542, 281.0981, 281.1418, 281.1855, 281.2295, 281.2732, 
    281.3169, 281.3787, 281.4487, 281.5188, 281.5889, 281.6589, 281.729, 
    281.7991, 281.8691, 281.9392, 282.0093, 282.0791, 282.1492, 282.2192, 
    282.2893, 282.3083, 282.2959, 282.2825, 282.2676, 282.251, 282.2327, 
    282.2124, 282.3513, 282.353, 282.3545, 282.3557, 282.3569, 282.3579, 
    282.3586, 282.3491, 281.8079, 281.7468, 281.6953, 281.6506, 281.6121, 
    281.5784, 281.5483, 281.5217, 281.4978, 281.4763, 281.4568, 281.439, 
    281.4229, 281.4153, 281.4155, 281.4158, 281.416, 281.416, 281.4163, 
    281.4165, 281.4167, 281.417, 281.4172, 281.4175, 281.4177, 281.418, 
    281.418, 281.4136, 281.4028, 281.3923, 281.3816, 281.3711, 281.3604, 
    281.3499, 281.3391, 281.3286, 281.3179, 281.3074, 281.2966, 281.2861, 
    281.2754, 281.2627, 281.2461, 281.2295, 281.2131, 281.1965, 281.1799, 
    281.1636, 281.147, 281.1304, 281.114, 281.0974, 281.0808, 281.0645, 
    281.0479, 281.0254, 280.9897, 280.9539, 280.9182, 280.8826, 280.8469, 
    280.8113, 280.7756, 280.74, 280.7043, 280.6687, 280.6331, 280.5972, 
    280.5615, 280.5254, 280.4878, 280.45, 280.4121, 280.3745, 280.3367, 
    280.2988, 280.2612, 280.2234, 280.1855, 280.1479, 280.1101, 280.0725, 
    280.0347, 279.9958, 279.9531, 279.9104, 279.8677, 279.8247, 279.782, 
    279.7393, 279.6965, 279.6538, 279.6108, 279.5681, 279.5254, 279.4827, 
    279.4397, 279.3928, 279.3169, 279.2407, 279.1648, 279.0889, 279.0127, 
    278.9368, 278.8608, 278.7847, 278.7087, 278.6328, 278.5566, 278.4807, 
    278.4045, 278.3325, 278.3198, 278.3071, 278.2944, 278.2817, 278.269, 
    278.2563, 278.2437, 278.231, 278.2183, 278.2056, 278.1926, 278.1799, 
    278.1672, 278.1545, 278.1807, 278.207, 278.2332, 278.2593, 278.2854, 
    278.3118, 278.3379, 278.364, 278.3901, 278.4163, 278.4426, 278.4688, 
    278.4949, 278.521, 278.5444, 278.5676, 278.5908, 278.6143, 278.6375, 
    278.6606, 278.6838, 278.707, 278.7302, 278.7537, 278.7769,
  276.197, 276.2397, 276.2827, 276.3254, 276.3684, 276.4111, 276.4541, 
    276.5039, 276.6018, 276.7, 276.7979, 276.896, 276.9939, 277.092, 
    277.1899, 277.2881, 277.386, 277.4841, 277.582, 277.6802, 277.7781, 
    277.8745, 277.9448, 278.0151, 278.0857, 278.156, 278.2263, 278.2966, 
    278.3669, 278.4375, 278.5078, 278.5781, 278.6484, 278.7188, 278.7893, 
    278.8596, 278.7297, 278.5999, 278.47, 278.3401, 278.21, 278.0801, 
    277.9502, 277.8203, 277.6904, 277.5605, 277.4307, 277.3008, 277.1709, 
    277.041, 277.1233, 277.2197, 277.3162, 277.4126, 277.509, 277.6055, 
    277.7019, 277.7983, 277.8948, 277.9912, 278.0876, 278.1841, 278.2805, 
    278.377, 278.5078, 278.6433, 278.7791, 278.9146, 279.0503, 279.1858, 
    279.3215, 279.457, 279.5928, 279.7285, 279.864, 279.9998, 280.1353, 
    280.271, 280.3247, 280.3599, 280.3948, 280.4299, 280.4648, 280.4998, 
    280.5349, 280.5698, 280.605, 280.6399, 280.6748, 280.71, 280.7449, 
    280.78, 280.8188, 280.8591, 280.8992, 280.9395, 280.9797, 281.02, 
    281.0601, 281.1003, 281.1406, 281.1809, 281.2209, 281.2612, 281.3015, 
    281.3418, 281.3948, 281.4536, 281.5125, 281.5715, 281.6304, 281.6892, 
    281.748, 281.8071, 281.866, 281.9248, 281.9836, 282.0427, 282.1016, 
    282.1604, 282.1741, 282.1599, 282.1445, 282.1279, 282.1101, 282.0908, 
    282.0698, 282.2917, 282.2976, 282.3027, 282.3071, 282.311, 282.3147, 
    282.3179, 282.3076, 281.739, 281.6907, 281.6475, 281.6084, 281.5732, 
    281.5413, 281.5122, 281.4854, 281.4607, 281.438, 281.417, 281.3975, 
    281.3794, 281.3687, 281.3645, 281.3606, 281.3564, 281.3523, 281.3484, 
    281.3442, 281.3401, 281.3362, 281.332, 281.3279, 281.324, 281.3198, 
    281.3157, 281.3125, 281.3103, 281.3081, 281.3059, 281.3035, 281.3013, 
    281.2991, 281.2969, 281.2947, 281.2925, 281.2903, 281.2881, 281.2859, 
    281.2837, 281.2788, 281.2695, 281.2605, 281.2512, 281.2422, 281.2329, 
    281.2239, 281.2146, 281.2056, 281.1963, 281.1873, 281.178, 281.1689, 
    281.1597, 281.1394, 281.095, 281.0503, 281.0056, 280.9609, 280.9165, 
    280.8718, 280.8271, 280.7825, 280.738, 280.6934, 280.6487, 280.604, 
    280.5593, 280.5168, 280.4797, 280.4429, 280.406, 280.3691, 280.3323, 
    280.2954, 280.2585, 280.2214, 280.1846, 280.1477, 280.1108, 280.074, 
    280.0371, 279.9993, 279.9585, 279.9175, 279.8767, 279.8359, 279.7949, 
    279.7542, 279.7131, 279.6724, 279.6313, 279.5906, 279.5496, 279.5088, 
    279.4678, 279.4231, 279.3503, 279.2776, 279.2048, 279.1323, 279.0596, 
    278.9868, 278.9141, 278.8416, 278.7688, 278.696, 278.6233, 278.5505, 
    278.478, 278.4087, 278.3921, 278.3752, 278.3586, 278.342, 278.3252, 
    278.3086, 278.2917, 278.2751, 278.2583, 278.2417, 278.2251, 278.2083, 
    278.1917, 278.1748, 278.1985, 278.2222, 278.2458, 278.2693, 278.293, 
    278.3167, 278.3403, 278.3638, 278.3875, 278.4111, 278.4348, 278.4585, 
    278.4819, 278.5056, 278.5203, 278.5342, 278.5481, 278.5623, 278.5762, 
    278.5901, 278.6042, 278.6182, 278.6321, 278.646, 278.6602,
  276.3877, 276.4355, 276.4834, 276.5312, 276.5789, 276.6267, 276.6746, 
    276.7288, 276.8286, 276.9282, 277.0278, 277.1277, 277.2273, 277.3269, 
    277.4268, 277.5264, 277.626, 277.7258, 277.8254, 277.925, 278.0247, 
    278.124, 278.218, 278.3123, 278.4062, 278.5002, 278.5942, 278.6882, 
    278.7822, 278.8762, 278.9702, 279.0642, 279.1582, 279.2524, 279.3464, 
    279.4404, 279.2761, 279.1121, 278.948, 278.7837, 278.6196, 278.4556, 
    278.2913, 278.1272, 277.9631, 277.7988, 277.6348, 277.4707, 277.3064, 
    277.1423, 277.21, 277.293, 277.376, 277.459, 277.542, 277.625, 277.708, 
    277.791, 277.874, 277.957, 278.04, 278.123, 278.2061, 278.2891, 278.4233, 
    278.5647, 278.7063, 278.8479, 278.9895, 279.1311, 279.2727, 279.4143, 
    279.5559, 279.6975, 279.8391, 279.9807, 280.1223, 280.2639, 280.3235, 
    280.3643, 280.4048, 280.4456, 280.4861, 280.5269, 280.5676, 280.6082, 
    280.6489, 280.6895, 280.7302, 280.7708, 280.8115, 280.8521, 280.8899, 
    280.9265, 280.9631, 280.9998, 281.0364, 281.073, 281.1099, 281.1465, 
    281.1831, 281.2197, 281.2563, 281.293, 281.3298, 281.3665, 281.4106, 
    281.4585, 281.5061, 281.554, 281.6018, 281.6494, 281.6973, 281.7449, 
    281.7927, 281.8406, 281.8882, 281.936, 281.9836, 282.0315, 282.0413, 
    282.0273, 282.0129, 281.9976, 281.9812, 281.9641, 281.9458, 282.2139, 
    282.2239, 282.2329, 282.241, 282.2483, 282.2546, 282.2605, 282.2493, 
    281.6909, 281.6494, 281.6108, 281.5747, 281.5413, 281.5098, 281.4805, 
    281.4529, 281.4268, 281.4021, 281.3789, 281.3569, 281.3362, 281.322, 
    281.3137, 281.3054, 281.2969, 281.2886, 281.2803, 281.272, 281.2634, 
    281.2551, 281.2468, 281.2385, 281.23, 281.2217, 281.2134, 281.2114, 
    281.2175, 281.2236, 281.23, 281.2361, 281.2422, 281.2485, 281.2546, 
    281.2607, 281.2671, 281.2732, 281.2793, 281.2854, 281.2917, 281.2949, 
    281.293, 281.2913, 281.2896, 281.2878, 281.2859, 281.2842, 281.2825, 
    281.2805, 281.2788, 281.2771, 281.2751, 281.2734, 281.2717, 281.2537, 
    281.2002, 281.1465, 281.093, 281.0393, 280.9858, 280.9324, 280.8787, 
    280.8252, 280.7715, 280.718, 280.6643, 280.6108, 280.5574, 280.5081, 
    280.4719, 280.436, 280.3999, 280.3638, 280.3279, 280.2917, 280.2556, 
    280.2197, 280.1836, 280.1475, 280.1116, 280.0754, 280.0393, 280.0027, 
    279.9639, 279.9248, 279.8857, 279.8469, 279.8079, 279.7688, 279.7297, 
    279.6909, 279.6519, 279.6128, 279.574, 279.5349, 279.4958, 279.4531, 
    279.3838, 279.3145, 279.2451, 279.1755, 279.1062, 279.0369, 278.9675, 
    278.8982, 278.8289, 278.7593, 278.6899, 278.6206, 278.5513, 278.4849, 
    278.4644, 278.4436, 278.4229, 278.4021, 278.3813, 278.3608, 278.3401, 
    278.3193, 278.2986, 278.2781, 278.2573, 278.2366, 278.2158, 278.1951, 
    278.2163, 278.2373, 278.2583, 278.2795, 278.3005, 278.3215, 278.3428, 
    278.3638, 278.3848, 278.406, 278.427, 278.448, 278.4692, 278.4902, 
    278.4961, 278.5007, 278.5054, 278.5103, 278.5149, 278.5198, 278.5244, 
    278.5291, 278.5339, 278.5386, 278.5435,
  276.5786, 276.6313, 276.6841, 276.7368, 276.7896, 276.8423, 276.895, 
    276.9539, 277.0552, 277.1565, 277.2578, 277.3591, 277.4607, 277.562, 
    277.6633, 277.7646, 277.866, 277.9673, 278.0686, 278.1699, 278.2715, 
    278.3738, 278.4915, 278.6091, 278.7268, 278.8445, 278.9622, 279.0798, 
    279.1975, 279.3152, 279.4329, 279.5505, 279.6682, 279.7859, 279.9036, 
    280.0212, 279.8228, 279.6243, 279.426, 279.2275, 279.0293, 278.8308, 
    278.6323, 278.4341, 278.2356, 278.0371, 277.8389, 277.6404, 277.4421, 
    277.2437, 277.2964, 277.366, 277.4355, 277.5051, 277.5747, 277.6443, 
    277.7139, 277.7834, 277.853, 277.9226, 277.9922, 278.0618, 278.1313, 
    278.2009, 278.3386, 278.4863, 278.6338, 278.7812, 278.929, 279.0764, 
    279.2241, 279.3716, 279.5193, 279.6667, 279.8142, 279.9619, 280.1094, 
    280.2571, 280.3223, 280.3687, 280.415, 280.4612, 280.5076, 280.554, 
    280.6001, 280.6465, 280.6929, 280.739, 280.7854, 280.8318, 280.8782, 
    280.9243, 280.9607, 280.9939, 281.0271, 281.0601, 281.0933, 281.1262, 
    281.1594, 281.1926, 281.2256, 281.2588, 281.2917, 281.325, 281.3582, 
    281.3911, 281.4268, 281.4634, 281.4998, 281.5364, 281.573, 281.6096, 
    281.6462, 281.6829, 281.7195, 281.7561, 281.7927, 281.8293, 281.866, 
    281.9026, 281.9097, 281.8987, 281.8872, 281.8752, 281.8628, 281.8501, 
    281.8367, 282.1072, 282.1213, 282.134, 282.1458, 282.1562, 282.166, 
    282.1748, 282.1624, 281.6553, 281.6177, 281.5818, 281.5474, 281.5144, 
    281.4829, 281.4526, 281.4233, 281.3955, 281.3684, 281.3425, 281.3176, 
    281.2935, 281.2754, 281.2627, 281.2502, 281.2375, 281.2249, 281.2122, 
    281.1995, 281.187, 281.1743, 281.1616, 281.1489, 281.1362, 281.1238, 
    281.1111, 281.1104, 281.1248, 281.1394, 281.1541, 281.1687, 281.1831, 
    281.1978, 281.2124, 281.2268, 281.2415, 281.2561, 281.2705, 281.2852, 
    281.2998, 281.311, 281.3167, 281.322, 281.3276, 281.3333, 281.3389, 
    281.3445, 281.3501, 281.3557, 281.3613, 281.3669, 281.3723, 281.3779, 
    281.3835, 281.3679, 281.3054, 281.2429, 281.1804, 281.1177, 281.0552, 
    280.9927, 280.9302, 280.8677, 280.8052, 280.7427, 280.6802, 280.6177, 
    280.5552, 280.4993, 280.4641, 280.429, 280.3938, 280.3586, 280.3235, 
    280.2881, 280.2529, 280.2178, 280.1826, 280.1475, 280.1121, 280.0769, 
    280.0417, 280.0061, 279.969, 279.9319, 279.895, 279.8579, 279.8208, 
    279.7837, 279.7466, 279.7095, 279.6724, 279.6353, 279.5981, 279.561, 
    279.5239, 279.4834, 279.4172, 279.3511, 279.2852, 279.219, 279.1531, 
    279.0869, 279.021, 278.9548, 278.8887, 278.8228, 278.7566, 278.6907, 
    278.6245, 278.561, 278.5364, 278.5117, 278.4871, 278.4624, 278.4377, 
    278.4131, 278.3882, 278.3635, 278.3389, 278.3142, 278.2896, 278.2649, 
    278.2402, 278.2156, 278.2339, 278.2524, 278.271, 278.2896, 278.3081, 
    278.3267, 278.3452, 278.3638, 278.3821, 278.4006, 278.4192, 278.4377, 
    278.4563, 278.4749, 278.4717, 278.4673, 278.4626, 278.4583, 278.4536, 
    278.4492, 278.4446, 278.4402, 278.4358, 278.4312, 278.4268,
  276.7695, 276.8271, 276.8848, 276.9424, 277.0002, 277.0579, 277.1155, 
    277.179, 277.282, 277.385, 277.4878, 277.5908, 277.6938, 277.7969, 
    277.8999, 278.0029, 278.106, 278.209, 278.312, 278.415, 278.5181, 
    278.6233, 278.7646, 278.906, 279.0474, 279.1887, 279.3301, 279.4714, 
    279.6125, 279.7539, 279.8953, 280.0366, 280.178, 280.3193, 280.4607, 
    280.6021, 280.3694, 280.1367, 279.9041, 279.6714, 279.4387, 279.2061, 
    278.9734, 278.7407, 278.5083, 278.2756, 278.043, 277.8103, 277.5776, 
    277.345, 277.3831, 277.4392, 277.4954, 277.5515, 277.6077, 277.6638, 
    277.72, 277.7761, 277.832, 277.8882, 277.9443, 278.0005, 278.0566, 
    278.1128, 278.2542, 278.4077, 278.5613, 278.7148, 278.8682, 279.0217, 
    279.1753, 279.3289, 279.4824, 279.636, 279.7896, 279.9429, 280.0964, 
    280.25, 280.321, 280.373, 280.425, 280.4771, 280.5288, 280.5808, 
    280.6328, 280.6848, 280.7368, 280.7888, 280.8408, 280.8926, 280.9446, 
    280.9966, 281.0317, 281.0613, 281.0908, 281.1204, 281.1499, 281.1794, 
    281.209, 281.2385, 281.2681, 281.2976, 281.3271, 281.3567, 281.3862, 
    281.4158, 281.4426, 281.468, 281.4937, 281.519, 281.5444, 281.5698, 
    281.5955, 281.6208, 281.6462, 281.6719, 281.6973, 281.7227, 281.748, 
    281.7737, 281.7793, 281.7732, 281.7668, 281.7605, 281.7539, 281.7471, 
    281.7402, 281.9524, 281.968, 281.9824, 281.9961, 282.009, 282.021, 
    282.0325, 282.0178, 281.6279, 281.5928, 281.5583, 281.5247, 281.4917, 
    281.4595, 281.4277, 281.3967, 281.3665, 281.3367, 281.3076, 281.2791, 
    281.2512, 281.2288, 281.2119, 281.1951, 281.178, 281.1611, 281.144, 
    281.1272, 281.1104, 281.0933, 281.0764, 281.0596, 281.0425, 281.0256, 
    281.0088, 281.0093, 281.0322, 281.0552, 281.0781, 281.1011, 281.124, 
    281.147, 281.1699, 281.1929, 281.2161, 281.239, 281.262, 281.2849, 
    281.3079, 281.3271, 281.3401, 281.353, 281.366, 281.3789, 281.3918, 
    281.4048, 281.4177, 281.4307, 281.4436, 281.4565, 281.4695, 281.4827, 
    281.4956, 281.4822, 281.4106, 281.3391, 281.2676, 281.1963, 281.1248, 
    281.0532, 280.9817, 280.9102, 280.8389, 280.7673, 280.6958, 280.6243, 
    280.553, 280.4907, 280.4563, 280.4219, 280.3877, 280.3533, 280.3188, 
    280.2847, 280.2502, 280.2158, 280.1816, 280.1472, 280.1128, 280.0784, 
    280.0442, 280.0095, 279.9744, 279.9392, 279.9041, 279.8689, 279.8337, 
    279.7983, 279.7632, 279.728, 279.6929, 279.6577, 279.6226, 279.5872, 
    279.552, 279.5134, 279.4507, 279.3879, 279.3252, 279.2625, 279.1997, 
    279.137, 279.0742, 279.0115, 278.9487, 278.886, 278.8232, 278.7605, 
    278.698, 278.6372, 278.6086, 278.5798, 278.5513, 278.5225, 278.4939, 
    278.4651, 278.4365, 278.4077, 278.3792, 278.3506, 278.3218, 278.2932, 
    278.2644, 278.2358, 278.2517, 278.2678, 278.2837, 278.2996, 278.3157, 
    278.3315, 278.3477, 278.3635, 278.3796, 278.3955, 278.4114, 278.4275, 
    278.4434, 278.4595, 278.4475, 278.4338, 278.4199, 278.4062, 278.3926, 
    278.3787, 278.365, 278.3513, 278.3374, 278.3237, 278.3101,
  276.9602, 277.0229, 277.0854, 277.1482, 277.2107, 277.2734, 277.3359, 
    277.4038, 277.5085, 277.6133, 277.7178, 277.8225, 277.9272, 278.032, 
    278.1365, 278.2412, 278.3459, 278.4507, 278.5552, 278.6599, 278.7646, 
    278.873, 279.0381, 279.2029, 279.3679, 279.533, 279.698, 279.8628, 
    280.0278, 280.1929, 280.3579, 280.5227, 280.6877, 280.8528, 281.0178, 
    281.1826, 280.9158, 280.6489, 280.3821, 280.1152, 279.8484, 279.5813, 
    279.3145, 279.0476, 278.7808, 278.5139, 278.2471, 277.9802, 277.7131, 
    277.4463, 277.4697, 277.5125, 277.5552, 277.5977, 277.6404, 277.6831, 
    277.7258, 277.7686, 277.8113, 277.854, 277.8967, 277.9392, 277.9819, 
    278.0247, 278.1697, 278.3291, 278.4885, 278.6482, 278.8076, 278.967, 
    279.1267, 279.2861, 279.4456, 279.605, 279.7646, 279.9241, 280.0835, 
    280.2432, 280.3198, 280.3774, 280.4351, 280.4927, 280.5503, 280.6079, 
    280.6655, 280.7231, 280.7808, 280.8384, 280.896, 280.9536, 281.0112, 
    281.0688, 281.1028, 281.1287, 281.1548, 281.1807, 281.2068, 281.2327, 
    281.2585, 281.2847, 281.3105, 281.3367, 281.3625, 281.3887, 281.4146, 
    281.4407, 281.4585, 281.4729, 281.4873, 281.5015, 281.5159, 281.5303, 
    281.5444, 281.5588, 281.573, 281.5874, 281.6018, 281.616, 281.6304, 
    281.6448, 281.6504, 281.6511, 281.6516, 281.6523, 281.6531, 281.6536, 
    281.6543, 281.6548, 281.6555, 281.6562, 281.6567, 281.6575, 281.6582, 
    281.6587, 281.6399, 281.6062, 281.5725, 281.5388, 281.5054, 281.4722, 
    281.4387, 281.4058, 281.3726, 281.3396, 281.3069, 281.2742, 281.2415, 
    281.209, 281.1821, 281.1609, 281.1399, 281.1187, 281.0974, 281.0762, 
    281.0549, 281.0337, 281.0125, 280.9912, 280.97, 280.9487, 280.9275, 
    280.9062, 280.9082, 280.9395, 280.9709, 281.0022, 281.0337, 281.0649, 
    281.0964, 281.1277, 281.1592, 281.1904, 281.2219, 281.2532, 281.2847, 
    281.3159, 281.3433, 281.3635, 281.3838, 281.4041, 281.4246, 281.4448, 
    281.4651, 281.4854, 281.5059, 281.5261, 281.5464, 281.5669, 281.5872, 
    281.6074, 281.5962, 281.5159, 281.4353, 281.355, 281.2747, 281.1941, 
    281.1138, 281.0332, 280.9529, 280.8723, 280.792, 280.7117, 280.6311, 
    280.5508, 280.4819, 280.4485, 280.415, 280.3816, 280.3479, 280.3145, 
    280.281, 280.2476, 280.2141, 280.1804, 280.147, 280.1135, 280.0801, 
    280.0464, 280.0129, 279.9797, 279.9465, 279.9131, 279.8799, 279.8464, 
    279.8132, 279.78, 279.7466, 279.7134, 279.6799, 279.6467, 279.6135, 
    279.5801, 279.5437, 279.4841, 279.4248, 279.3652, 279.3059, 279.2466, 
    279.187, 279.1277, 279.0684, 279.0088, 278.9495, 278.8901, 278.8306, 
    278.7712, 278.7134, 278.6807, 278.6482, 278.6155, 278.5828, 278.55, 
    278.5173, 278.4846, 278.4521, 278.4194, 278.3867, 278.354, 278.3213, 
    278.2888, 278.2561, 278.2695, 278.283, 278.2964, 278.3098, 278.3232, 
    278.3367, 278.3501, 278.3635, 278.377, 278.3904, 278.4038, 278.4172, 
    278.4307, 278.4441, 278.4233, 278.4004, 278.3772, 278.3542, 278.3313, 
    278.3083, 278.2852, 278.2622, 278.2393, 278.2163, 278.1931,
  276.9517, 277.0115, 277.0713, 277.1311, 277.1909, 277.2507, 277.3105, 
    277.3748, 277.4697, 277.5647, 277.6594, 277.7544, 277.8491, 277.9441, 
    278.0388, 278.1338, 278.2285, 278.3235, 278.4182, 278.5132, 278.6079, 
    278.707, 278.8667, 279.0266, 279.1865, 279.3462, 279.5061, 279.666, 
    279.8257, 279.9856, 280.1455, 280.3052, 280.4651, 280.625, 280.7847, 
    280.9446, 280.7073, 280.47, 280.2324, 279.9951, 279.7578, 279.5205, 
    279.283, 279.0457, 278.8083, 278.571, 278.3335, 278.0962, 277.8589, 
    277.6216, 277.6443, 277.6843, 277.7246, 277.7646, 277.8049, 277.845, 
    277.885, 277.9253, 277.9653, 278.0056, 278.0457, 278.0859, 278.126, 
    278.166, 278.304, 278.4556, 278.6074, 278.759, 278.9109, 279.0625, 
    279.2141, 279.366, 279.5176, 279.6694, 279.821, 279.9729, 280.1245, 
    280.2764, 280.356, 280.4189, 280.4819, 280.5449, 280.6079, 280.6709, 
    280.7339, 280.7969, 280.8599, 280.9229, 280.9858, 281.0488, 281.1118, 
    281.1748, 281.21, 281.2356, 281.2615, 281.2871, 281.3127, 281.3386, 
    281.3643, 281.3899, 281.4158, 281.4414, 281.467, 281.4929, 281.5186, 
    281.5442, 281.5508, 281.5488, 281.5466, 281.5444, 281.5425, 281.5403, 
    281.5381, 281.5361, 281.5339, 281.5317, 281.5298, 281.5276, 281.5254, 
    281.5232, 281.5217, 281.5203, 281.519, 281.5176, 281.5164, 281.5149, 
    281.5137, 281.5122, 281.511, 281.5095, 281.5083, 281.5068, 281.5056, 
    281.5042, 281.4902, 281.4663, 281.4426, 281.4187, 281.395, 281.3713, 
    281.3474, 281.3237, 281.2998, 281.2761, 281.2522, 281.2285, 281.2048, 
    281.1809, 281.1599, 281.1414, 281.1228, 281.1042, 281.0859, 281.0674, 
    281.0488, 281.0305, 281.012, 280.9934, 280.9751, 280.9565, 280.938, 
    280.9194, 280.9236, 280.9565, 280.9897, 281.0227, 281.0557, 281.0886, 
    281.1218, 281.1548, 281.1877, 281.2207, 281.2539, 281.2869, 281.3198, 
    281.353, 281.3813, 281.4019, 281.4224, 281.4429, 281.4634, 281.4839, 
    281.5044, 281.5249, 281.5454, 281.5659, 281.5864, 281.6069, 281.6274, 
    281.6482, 281.6355, 281.5498, 281.4641, 281.3784, 281.2927, 281.207, 
    281.1213, 281.0356, 280.95, 280.8643, 280.7786, 280.6929, 280.6072, 
    280.5215, 280.4492, 280.4167, 280.3843, 280.3518, 280.3193, 280.2869, 
    280.2544, 280.2219, 280.1895, 280.157, 280.1245, 280.092, 280.0596, 
    280.0271, 279.9958, 279.969, 279.9421, 279.9153, 279.8884, 279.8616, 
    279.8347, 279.8081, 279.7812, 279.7544, 279.7275, 279.7007, 279.6738, 
    279.647, 279.6162, 279.5562, 279.4961, 279.436, 279.376, 279.3159, 
    279.2559, 279.1958, 279.136, 279.0759, 279.0159, 278.9558, 278.8958, 
    278.8357, 278.7773, 278.7415, 278.7058, 278.6699, 278.6343, 278.5986, 
    278.5627, 278.5271, 278.4915, 278.4556, 278.4199, 278.3843, 278.3484, 
    278.3127, 278.2771, 278.2893, 278.3015, 278.314, 278.3262, 278.3384, 
    278.3508, 278.363, 278.3755, 278.3877, 278.3999, 278.4124, 278.4246, 
    278.437, 278.4492, 278.4343, 278.4177, 278.4011, 278.3845, 278.3679, 
    278.3513, 278.3347, 278.3181, 278.3015, 278.2849, 278.2683,
  276.8931, 276.948, 277.0032, 277.0583, 277.1135, 277.1685, 277.2236, 
    277.2822, 277.3643, 277.4465, 277.5286, 277.6108, 277.6929, 277.7751, 
    277.8574, 277.9395, 278.0217, 278.1038, 278.186, 278.2681, 278.3503, 
    278.4365, 278.584, 278.7314, 278.8789, 279.0264, 279.1738, 279.3213, 
    279.4688, 279.6162, 279.7637, 279.9111, 280.0586, 280.2061, 280.3535, 
    280.501, 280.3093, 280.1174, 279.9255, 279.7336, 279.5417, 279.3499, 
    279.158, 278.9663, 278.7744, 278.5825, 278.3906, 278.1987, 278.0068, 
    277.8152, 277.8408, 277.8811, 277.9216, 277.9619, 278.0022, 278.0425, 
    278.0828, 278.123, 278.1636, 278.2039, 278.2441, 278.2844, 278.3247, 
    278.365, 278.4929, 278.6335, 278.7739, 278.9146, 279.0549, 279.1956, 
    279.3359, 279.4766, 279.6169, 279.7576, 279.8979, 280.0386, 280.179, 
    280.3196, 280.4014, 280.4697, 280.5381, 280.6062, 280.6746, 280.7429, 
    280.8113, 280.8796, 280.9478, 281.0161, 281.0845, 281.1528, 281.2212, 
    281.2896, 281.3262, 281.3525, 281.3787, 281.405, 281.4314, 281.4575, 
    281.4839, 281.5103, 281.5364, 281.5627, 281.5889, 281.6152, 281.6416, 
    281.6677, 281.6624, 281.6423, 281.6226, 281.6025, 281.5828, 281.563, 
    281.543, 281.5232, 281.5032, 281.4834, 281.4634, 281.4436, 281.4236, 
    281.4038, 281.3928, 281.387, 281.3811, 281.3752, 281.3694, 281.3638, 
    281.3579, 281.3521, 281.3462, 281.3403, 281.3345, 281.3289, 281.323, 
    281.3171, 281.3081, 281.2964, 281.2847, 281.2729, 281.2612, 281.2498, 
    281.238, 281.2263, 281.2146, 281.2029, 281.1914, 281.1797, 281.168, 
    281.1562, 281.1436, 281.1294, 281.1155, 281.1016, 281.0876, 281.0735, 
    281.0596, 281.0457, 281.0317, 281.0176, 281.0037, 280.9897, 280.9758, 
    280.9617, 280.9683, 281.0012, 281.0342, 281.0674, 281.1003, 281.1333, 
    281.1663, 281.1992, 281.2322, 281.2651, 281.2981, 281.3311, 281.364, 
    281.3972, 281.4248, 281.4438, 281.4626, 281.4817, 281.5005, 281.5195, 
    281.5383, 281.5574, 281.5762, 281.5952, 281.614, 281.6331, 281.6519, 
    281.6709, 281.6558, 281.5657, 281.4758, 281.3857, 281.2957, 281.2058, 
    281.1157, 281.0256, 280.9355, 280.8457, 280.7556, 280.6655, 280.5757, 
    280.4856, 280.4102, 280.3789, 280.3474, 280.3162, 280.2847, 280.2534, 
    280.2219, 280.1907, 280.1592, 280.1279, 280.0964, 280.0652, 280.0337, 
    280.0024, 279.9731, 279.9541, 279.9348, 279.9158, 279.8965, 279.8772, 
    279.8582, 279.8389, 279.8198, 279.8005, 279.7812, 279.7622, 279.7429, 
    279.7239, 279.6992, 279.6377, 279.5759, 279.5144, 279.4529, 279.3911, 
    279.3296, 279.2678, 279.2063, 279.1445, 279.083, 279.0212, 278.9597, 
    278.8982, 278.8379, 278.7993, 278.7607, 278.7222, 278.6836, 278.645, 
    278.6064, 278.5681, 278.5295, 278.491, 278.4524, 278.4138, 278.3752, 
    278.3367, 278.2981, 278.3096, 278.321, 278.3328, 278.3442, 278.3557, 
    278.3672, 278.3789, 278.3904, 278.4019, 278.4133, 278.425, 278.4365, 
    278.448, 278.4595, 278.4543, 278.448, 278.4417, 278.4355, 278.4292, 
    278.4229, 278.4165, 278.4102, 278.4041, 278.3977, 278.3914,
  276.8342, 276.8848, 276.9351, 276.9854, 277.0359, 277.0862, 277.1367, 
    277.1895, 277.2588, 277.3284, 277.3979, 277.4673, 277.5369, 277.6062, 
    277.6758, 277.7454, 277.8147, 277.8843, 277.9536, 278.0232, 278.0928, 
    278.1663, 278.3013, 278.4365, 278.5715, 278.7065, 278.8418, 278.9768, 
    279.1118, 279.2471, 279.3821, 279.5171, 279.6523, 279.7874, 279.9224, 
    280.0576, 279.9111, 279.7649, 279.6184, 279.4722, 279.3259, 279.1794, 
    279.0332, 278.8867, 278.7405, 278.594, 278.4478, 278.3015, 278.155, 
    278.0088, 278.0376, 278.0781, 278.1184, 278.1589, 278.1995, 278.24, 
    278.2805, 278.321, 278.3616, 278.4021, 278.4426, 278.4829, 278.5234, 
    278.564, 278.6821, 278.8115, 278.9407, 279.0701, 279.1992, 279.3286, 
    279.4578, 279.5872, 279.7163, 279.8457, 279.9749, 280.1042, 280.2334, 
    280.3628, 280.4468, 280.5205, 280.594, 280.6677, 280.7412, 280.8149, 
    280.8887, 280.9622, 281.0359, 281.1094, 281.1831, 281.2568, 281.3303, 
    281.4041, 281.4426, 281.4692, 281.4961, 281.5229, 281.5498, 281.5767, 
    281.6035, 281.6304, 281.6572, 281.6838, 281.7107, 281.7375, 281.7644, 
    281.7913, 281.7737, 281.7361, 281.6985, 281.6609, 281.623, 281.5854, 
    281.5479, 281.5103, 281.4727, 281.4348, 281.3972, 281.3596, 281.322, 
    281.2844, 281.2637, 281.2534, 281.2432, 281.2329, 281.2227, 281.2124, 
    281.2021, 281.1919, 281.1816, 281.1711, 281.1609, 281.1506, 281.1404, 
    281.1301, 281.126, 281.1262, 281.1267, 281.1272, 281.1277, 281.1282, 
    281.1284, 281.1289, 281.1294, 281.1299, 281.1304, 281.1306, 281.1311, 
    281.1316, 281.127, 281.1177, 281.1082, 281.0986, 281.0891, 281.0798, 
    281.0703, 281.0608, 281.0513, 281.0417, 281.0325, 281.0229, 281.0134, 
    281.0039, 281.0129, 281.0459, 281.0789, 281.1118, 281.1448, 281.1777, 
    281.2107, 281.2437, 281.2766, 281.3096, 281.3425, 281.3755, 281.4084, 
    281.4414, 281.4685, 281.4858, 281.5032, 281.5205, 281.5376, 281.5549, 
    281.5723, 281.5896, 281.6069, 281.6243, 281.6416, 281.6589, 281.6763, 
    281.6936, 281.676, 281.5818, 281.4873, 281.3931, 281.2988, 281.2043, 
    281.1101, 281.0156, 280.9214, 280.8271, 280.7327, 280.6384, 280.5439, 
    280.4497, 280.3713, 280.3411, 280.3108, 280.2805, 280.2502, 280.22, 
    280.1897, 280.1594, 280.1292, 280.0986, 280.0684, 280.0381, 280.0078, 
    279.9775, 279.9507, 279.9392, 279.9277, 279.916, 279.9045, 279.8931, 
    279.8813, 279.8699, 279.8584, 279.8467, 279.8352, 279.8235, 279.812, 
    279.8005, 279.7825, 279.7192, 279.656, 279.5928, 279.5295, 279.4663, 
    279.4031, 279.3398, 279.2766, 279.2134, 279.1501, 279.0869, 279.0237, 
    278.9604, 278.8987, 278.8572, 278.8159, 278.7744, 278.7332, 278.6917, 
    278.6504, 278.6089, 278.5676, 278.5261, 278.4849, 278.4434, 278.4021, 
    278.3606, 278.3193, 278.3301, 278.3408, 278.3516, 278.3623, 278.373, 
    278.3838, 278.3945, 278.4053, 278.416, 278.4268, 278.4375, 278.4482, 
    278.459, 278.47, 278.4744, 278.4783, 278.4824, 278.4863, 278.4902, 
    278.4944, 278.4983, 278.5024, 278.5063, 278.5105, 278.5144,
  276.7756, 276.8213, 276.8669, 276.9126, 276.9583, 277.0039, 277.0496, 
    277.0967, 277.1536, 277.2102, 277.2671, 277.324, 277.3806, 277.4375, 
    277.4941, 277.551, 277.6079, 277.6646, 277.7214, 277.7783, 277.835, 
    277.896, 278.0188, 278.1414, 278.2642, 278.387, 278.5095, 278.6323, 
    278.7551, 278.8777, 279.0005, 279.1233, 279.2458, 279.3687, 279.4915, 
    279.614, 279.5132, 279.4124, 279.3115, 279.2107, 279.1099, 279.009, 
    278.9082, 278.8074, 278.7065, 278.6057, 278.5049, 278.4041, 278.3032, 
    278.2024, 278.2341, 278.2749, 278.3154, 278.3562, 278.397, 278.4375, 
    278.4783, 278.5188, 278.5596, 278.6003, 278.6409, 278.6816, 278.7222, 
    278.7629, 278.8713, 278.9893, 279.1074, 279.2256, 279.3435, 279.4617, 
    279.5796, 279.6978, 279.8157, 279.9338, 280.0518, 280.1699, 280.2878, 
    280.406, 280.4922, 280.5713, 280.6501, 280.729, 280.8081, 280.887, 
    280.9658, 281.0449, 281.1238, 281.2026, 281.2817, 281.3606, 281.4397, 
    281.5186, 281.5588, 281.5862, 281.6135, 281.6409, 281.6682, 281.6958, 
    281.7231, 281.7505, 281.7778, 281.8052, 281.8325, 281.8601, 281.8875, 
    281.9148, 281.8853, 281.8298, 281.7744, 281.719, 281.6636, 281.6082, 
    281.5527, 281.4973, 281.4419, 281.3865, 281.3311, 281.2756, 281.2202, 
    281.1648, 281.1348, 281.1201, 281.1052, 281.0906, 281.0759, 281.061, 
    281.0464, 281.0315, 281.0168, 281.0022, 280.9873, 280.9727, 280.9578, 
    280.9431, 280.9438, 280.9563, 280.9688, 280.9814, 280.9939, 281.0066, 
    281.019, 281.0315, 281.0442, 281.0566, 281.0693, 281.0818, 281.0942, 
    281.1069, 281.1106, 281.1057, 281.1008, 281.0957, 281.0908, 281.0859, 
    281.0808, 281.0759, 281.071, 281.0659, 281.061, 281.0562, 281.051, 
    281.0461, 281.0579, 281.0906, 281.1235, 281.1565, 281.1895, 281.2224, 
    281.2551, 281.2881, 281.321, 281.354, 281.3867, 281.4197, 281.4526, 
    281.4856, 281.512, 281.5278, 281.5435, 281.5591, 281.575, 281.5906, 
    281.6064, 281.6221, 281.6377, 281.6536, 281.6692, 281.6851, 281.7007, 
    281.7163, 281.6963, 281.5977, 281.499, 281.4004, 281.3018, 281.2031, 
    281.1045, 281.0056, 280.907, 280.8083, 280.7097, 280.6111, 280.5125, 
    280.4138, 280.3325, 280.3032, 280.2739, 280.2449, 280.2156, 280.1865, 
    280.1572, 280.1279, 280.0989, 280.0696, 280.0405, 280.0112, 279.9819, 
    279.9529, 279.9282, 279.9243, 279.9204, 279.9165, 279.9126, 279.9087, 
    279.9048, 279.9009, 279.8967, 279.8928, 279.8889, 279.885, 279.8811, 
    279.8772, 279.8657, 279.8008, 279.7358, 279.6711, 279.6062, 279.5415, 
    279.4766, 279.4119, 279.3469, 279.2822, 279.2173, 279.1526, 279.0876, 
    279.0227, 278.9592, 278.915, 278.8708, 278.8267, 278.7825, 278.7383, 
    278.6941, 278.6499, 278.6057, 278.5613, 278.5171, 278.4729, 278.4287, 
    278.3845, 278.3403, 278.3503, 278.3604, 278.3704, 278.3804, 278.3904, 
    278.4004, 278.4102, 278.4202, 278.4302, 278.4402, 278.4502, 278.4602, 
    278.4702, 278.4802, 278.4941, 278.5085, 278.5229, 278.5374, 278.5515, 
    278.5659, 278.5803, 278.5945, 278.6089, 278.6233, 278.6375,
  276.717, 276.7578, 276.7988, 276.8398, 276.8806, 276.9216, 276.9626, 
    277.0039, 277.0481, 277.092, 277.1362, 277.1804, 277.2246, 277.2686, 
    277.3127, 277.3569, 277.4009, 277.4451, 277.4893, 277.5332, 277.5774, 
    277.6257, 277.7361, 277.8464, 277.9568, 278.0671, 278.1775, 278.2878, 
    278.3982, 278.5085, 278.6189, 278.7292, 278.8396, 278.95, 279.0603, 
    279.1707, 279.1152, 279.0598, 279.0046, 278.9492, 278.8938, 278.8386, 
    278.7832, 278.728, 278.6726, 278.6172, 278.562, 278.5066, 278.4512, 
    278.396, 278.4309, 278.4717, 278.5125, 278.5535, 278.5942, 278.635, 
    278.676, 278.7168, 278.7576, 278.7986, 278.8394, 278.8801, 278.9211, 
    278.9619, 279.0605, 279.1672, 279.2742, 279.3809, 279.4878, 279.5945, 
    279.7014, 279.8083, 279.915, 280.022, 280.1287, 280.2356, 280.3423, 
    280.4492, 280.5376, 280.6218, 280.7063, 280.7905, 280.8748, 280.959, 
    281.0432, 281.1274, 281.2117, 281.2961, 281.3804, 281.4646, 281.5488, 
    281.6331, 281.675, 281.7031, 281.731, 281.7588, 281.7869, 281.8147, 
    281.8428, 281.8706, 281.8987, 281.9265, 281.9543, 281.9824, 282.0103, 
    282.0383, 281.9966, 281.9236, 281.8503, 281.7771, 281.7039, 281.6309, 
    281.5576, 281.4844, 281.4111, 281.3381, 281.2649, 281.1917, 281.1184, 
    281.0454, 281.0059, 280.9866, 280.9675, 280.9482, 280.929, 280.9099, 
    280.8906, 280.8713, 280.8521, 280.833, 280.8137, 280.7944, 280.7754, 
    280.7561, 280.7615, 280.7861, 280.8108, 280.8357, 280.8604, 280.885, 
    280.9097, 280.9343, 280.959, 280.9836, 281.0083, 281.033, 281.0576, 
    281.0823, 281.0942, 281.094, 281.0935, 281.093, 281.0925, 281.092, 
    281.0916, 281.0911, 281.0906, 281.0901, 281.0898, 281.0894, 281.0889, 
    281.0884, 281.1025, 281.1353, 281.1682, 281.2012, 281.2339, 281.2668, 
    281.2998, 281.3325, 281.3655, 281.3982, 281.4312, 281.4641, 281.4968, 
    281.5298, 281.5557, 281.5698, 281.5837, 281.5979, 281.6121, 281.6262, 
    281.6404, 281.6545, 281.6685, 281.6826, 281.6968, 281.7109, 281.7251, 
    281.7393, 281.7168, 281.6138, 281.5107, 281.4077, 281.3047, 281.2017, 
    281.0989, 280.9958, 280.8928, 280.7898, 280.6868, 280.5837, 280.4807, 
    280.3777, 280.2935, 280.2654, 280.2373, 280.2092, 280.1812, 280.1528, 
    280.1248, 280.0967, 280.0686, 280.0405, 280.0125, 279.9841, 279.9561, 
    279.928, 279.9058, 279.9097, 279.9133, 279.917, 279.9207, 279.9243, 
    279.928, 279.9316, 279.9353, 279.9392, 279.9429, 279.9465, 279.9502, 
    279.9539, 279.9487, 279.8823, 279.8159, 279.7495, 279.6831, 279.6167, 
    279.5503, 279.4836, 279.4172, 279.3508, 279.2844, 279.218, 279.1516, 
    279.0852, 279.02, 278.9729, 278.9258, 278.8789, 278.8318, 278.7847, 
    278.7378, 278.6907, 278.6436, 278.5967, 278.5496, 278.5027, 278.4556, 
    278.4084, 278.3616, 278.3706, 278.3799, 278.3892, 278.3984, 278.4075, 
    278.4167, 278.426, 278.4353, 278.4443, 278.4536, 278.4629, 278.4722, 
    278.4812, 278.4905, 278.5142, 278.5388, 278.5635, 278.5881, 278.6128, 
    278.6375, 278.6621, 278.6868, 278.7114, 278.7361, 278.7607,
  276.6582, 276.6946, 276.7307, 276.7668, 276.8032, 276.8394, 276.8755, 
    276.9111, 276.9426, 276.9741, 277.0054, 277.0369, 277.0684, 277.0999, 
    277.1311, 277.1626, 277.1941, 277.2253, 277.2568, 277.2883, 277.3198, 
    277.3552, 277.4534, 277.5513, 277.6492, 277.7473, 277.8452, 277.9431, 
    278.0413, 278.1392, 278.2371, 278.3352, 278.4331, 278.531, 278.6292, 
    278.7271, 278.7173, 278.7075, 278.6975, 278.6877, 278.678, 278.6682, 
    278.6582, 278.6484, 278.6387, 278.6289, 278.6191, 278.6091, 278.5994, 
    278.5896, 278.6274, 278.6685, 278.7095, 278.7505, 278.7915, 278.8325, 
    278.8735, 278.9146, 278.9556, 278.9968, 279.0378, 279.0789, 279.1199, 
    279.1609, 279.2495, 279.3452, 279.4409, 279.5364, 279.6321, 279.7275, 
    279.8232, 279.9187, 280.0144, 280.1101, 280.2056, 280.3013, 280.3967, 
    280.4924, 280.583, 280.6726, 280.7622, 280.8518, 280.9414, 281.031, 
    281.1206, 281.2102, 281.2998, 281.3894, 281.479, 281.5684, 281.658, 
    281.7476, 281.7915, 281.8198, 281.8484, 281.877, 281.9053, 281.9338, 
    281.9624, 281.9907, 282.0193, 282.0479, 282.0762, 282.1047, 282.1333, 
    282.1616, 282.1082, 282.0171, 281.9263, 281.8352, 281.7444, 281.6533, 
    281.5625, 281.4714, 281.3806, 281.2896, 281.1987, 281.1077, 281.0168, 
    280.9258, 280.877, 280.8533, 280.8296, 280.8059, 280.7822, 280.7585, 
    280.7349, 280.7112, 280.6875, 280.6638, 280.6401, 280.6165, 280.5928, 
    280.5691, 280.5793, 280.6162, 280.6531, 280.6897, 280.7266, 280.7634, 
    280.8, 280.8369, 280.8738, 280.9104, 280.9473, 280.9839, 281.0208, 
    281.0576, 281.0779, 281.082, 281.0862, 281.0901, 281.0942, 281.0981, 
    281.1023, 281.1062, 281.1104, 281.1145, 281.1184, 281.1226, 281.1265, 
    281.1306, 281.1472, 281.1799, 281.2129, 281.2456, 281.2786, 281.3113, 
    281.3442, 281.377, 281.4099, 281.4426, 281.4756, 281.5083, 281.541, 
    281.574, 281.5991, 281.6116, 281.6243, 281.6367, 281.6492, 281.6619, 
    281.6743, 281.6868, 281.6995, 281.7119, 281.7244, 281.7368, 281.7495, 
    281.762, 281.7371, 281.6296, 281.5225, 281.415, 281.3079, 281.2004, 
    281.093, 280.9858, 280.8784, 280.7712, 280.6638, 280.5564, 280.4492, 
    280.3418, 280.2546, 280.2275, 280.2007, 280.1736, 280.1465, 280.1194, 
    280.0925, 280.0654, 280.0383, 280.0112, 279.9844, 279.9573, 279.9302, 
    279.9033, 279.8833, 279.8948, 279.906, 279.9172, 279.9287, 279.9399, 
    279.9514, 279.9626, 279.9739, 279.9854, 279.9966, 280.0078, 280.0193, 
    280.0305, 280.032, 279.9639, 279.896, 279.8279, 279.7598, 279.6919, 
    279.6238, 279.5557, 279.4878, 279.4197, 279.3516, 279.2837, 279.2156, 
    279.1475, 279.0806, 279.0308, 278.981, 278.9312, 278.8811, 278.8313, 
    278.7815, 278.7317, 278.6816, 278.6318, 278.582, 278.5322, 278.4824, 
    278.4324, 278.3826, 278.3911, 278.3994, 278.408, 278.4163, 278.4248, 
    278.4333, 278.4417, 278.4502, 278.4585, 278.467, 278.4756, 278.4839, 
    278.4924, 278.5007, 278.5342, 278.5691, 278.604, 278.6389, 278.6741, 
    278.709, 278.7439, 278.7788, 278.8137, 278.8489, 278.8838,
  276.5996, 276.6311, 276.6626, 276.6941, 276.7256, 276.7571, 276.7886, 
    276.8184, 276.8372, 276.856, 276.8748, 276.8933, 276.9121, 276.9309, 
    276.9497, 276.9683, 276.9871, 277.0059, 277.0247, 277.0432, 277.062, 
    277.085, 277.1707, 277.2561, 277.3418, 277.4275, 277.5129, 277.5986, 
    277.6843, 277.7698, 277.8555, 277.9412, 278.0266, 278.1123, 278.198, 
    278.2834, 278.3193, 278.355, 278.3906, 278.4263, 278.4619, 278.4976, 
    278.5334, 278.5691, 278.6047, 278.6404, 278.676, 278.7119, 278.7476, 
    278.7832, 278.824, 278.8652, 278.9065, 278.9478, 278.989, 279.03, 
    279.0713, 279.1125, 279.1538, 279.1948, 279.2361, 279.2773, 279.3186, 
    279.3599, 279.4387, 279.5232, 279.6074, 279.6919, 279.7764, 279.8606, 
    279.9451, 280.0293, 280.1138, 280.1982, 280.2825, 280.3669, 280.4512, 
    280.5356, 280.6287, 280.7234, 280.8184, 280.9133, 281.0081, 281.103, 
    281.198, 281.2927, 281.3877, 281.4827, 281.5774, 281.6724, 281.7673, 
    281.8623, 281.9077, 281.9368, 281.9658, 281.9949, 282.0239, 282.053, 
    282.082, 282.1111, 282.1399, 282.1689, 282.198, 282.2271, 282.2561, 
    282.2852, 282.2195, 282.1108, 282.0022, 281.8933, 281.7847, 281.676, 
    281.5674, 281.4585, 281.3499, 281.2412, 281.1326, 281.0237, 280.915, 
    280.8064, 280.748, 280.7197, 280.6917, 280.6636, 280.6355, 280.6072, 
    280.5791, 280.551, 280.5227, 280.4946, 280.4666, 280.4385, 280.4102, 
    280.3821, 280.3972, 280.4463, 280.4951, 280.5439, 280.5928, 280.6418, 
    280.6907, 280.7395, 280.7883, 280.8374, 280.8862, 280.9351, 280.9839, 
    281.033, 281.0615, 281.0701, 281.0786, 281.0872, 281.0957, 281.1042, 
    281.113, 281.1216, 281.1301, 281.1387, 281.1472, 281.1558, 281.1643, 
    281.1729, 281.1919, 281.2246, 281.2576, 281.2903, 281.323, 281.356, 
    281.3887, 281.4214, 281.4543, 281.4871, 281.5198, 281.5525, 281.5854, 
    281.6182, 281.6428, 281.6536, 281.6646, 281.6755, 281.6865, 281.6973, 
    281.7083, 281.7192, 281.7302, 281.741, 281.752, 281.7629, 281.7739, 
    281.7847, 281.7573, 281.6458, 281.5342, 281.4224, 281.3108, 281.1992, 
    281.0874, 280.9758, 280.8643, 280.7524, 280.6409, 280.5293, 280.4175, 
    280.3059, 280.2158, 280.1897, 280.1638, 280.1379, 280.1121, 280.0859, 
    280.0601, 280.0342, 280.0081, 279.9822, 279.9563, 279.9304, 279.9043, 
    279.8784, 279.8608, 279.8799, 279.8989, 279.9177, 279.9368, 279.9556, 
    279.9746, 279.9937, 280.0125, 280.0315, 280.0503, 280.0693, 280.0884, 
    280.1072, 280.1152, 280.0454, 279.9758, 279.9062, 279.8367, 279.7668, 
    279.6973, 279.6277, 279.5581, 279.4885, 279.4187, 279.3491, 279.2795, 
    279.21, 279.1414, 279.0886, 279.0359, 278.9832, 278.9307, 278.8779, 
    278.8252, 278.7725, 278.7197, 278.6672, 278.6145, 278.5618, 278.509, 
    278.4563, 278.4038, 278.4114, 278.4189, 278.4268, 278.4343, 278.4421, 
    278.4497, 278.4575, 278.4651, 278.4729, 278.4805, 278.488, 278.4958, 
    278.5034, 278.5112, 278.5542, 278.5994, 278.6448, 278.6899, 278.7351, 
    278.7805, 278.8257, 278.8711, 278.9163, 278.9617, 279.0068,
  276.5581, 276.5813, 276.6064, 276.6357, 276.6648, 276.6941, 276.7231, 
    276.7507, 276.7668, 276.7832, 276.7993, 276.8154, 276.8315, 276.8479, 
    276.864, 276.8801, 276.8982, 276.9187, 276.939, 276.9595, 276.9797, 
    277.0039, 277.0837, 277.1638, 277.2439, 277.3237, 277.4038, 277.4836, 
    277.5637, 277.6436, 277.7227, 277.801, 277.8794, 277.9578, 278.0361, 
    278.1145, 278.1602, 278.2058, 278.2517, 278.2974, 278.343, 278.3887, 
    278.4346, 278.4802, 278.5325, 278.5881, 278.6436, 278.699, 278.7546, 
    278.8101, 278.8613, 278.9126, 278.9639, 279.0149, 279.0662, 279.1172, 
    279.1685, 279.2195, 279.2778, 279.3381, 279.3984, 279.4585, 279.5188, 
    279.5791, 279.6709, 279.7671, 279.8635, 279.9597, 280.0562, 280.1526, 
    280.2488, 280.3452, 280.4102, 280.4719, 280.5337, 280.5955, 280.6572, 
    280.719, 280.791, 280.8655, 280.9399, 281.0144, 281.0889, 281.1633, 
    281.2378, 281.3125, 281.4055, 281.4983, 281.5911, 281.6838, 281.7766, 
    281.8694, 281.9175, 281.9507, 281.9839, 282.0171, 282.0503, 282.0833, 
    282.1165, 282.1482, 282.1689, 282.1899, 282.2107, 282.2317, 282.2524, 
    282.2732, 282.2073, 282.1018, 281.9961, 281.8906, 281.7852, 281.6797, 
    281.574, 281.468, 281.3606, 281.2532, 281.1455, 281.0381, 280.9307, 
    280.823, 280.762, 280.729, 280.696, 280.6628, 280.6299, 280.5967, 
    280.5637, 280.5356, 280.5166, 280.4978, 280.4788, 280.46, 280.4409, 
    280.4221, 280.4436, 280.4966, 280.5498, 280.6028, 280.6558, 280.7087, 
    280.762, 280.8147, 280.8672, 280.9199, 280.9724, 281.0249, 281.0774, 
    281.1301, 281.1638, 281.179, 281.1941, 281.2092, 281.2241, 281.2393, 
    281.2544, 281.2651, 281.2727, 281.28, 281.2876, 281.2949, 281.3025, 
    281.3098, 281.3264, 281.3545, 281.3826, 281.4106, 281.4387, 281.4668, 
    281.4949, 281.5212, 281.5466, 281.572, 281.5974, 281.6228, 281.6482, 
    281.6738, 281.6917, 281.6973, 281.7029, 281.7087, 281.7144, 281.72, 
    281.7256, 281.7273, 281.728, 281.7288, 281.7295, 281.7302, 281.731, 
    281.7317, 281.6982, 281.5894, 281.4802, 281.3713, 281.2625, 281.1536, 
    281.0447, 280.9399, 280.8357, 280.7312, 280.627, 280.5227, 280.4185, 
    280.3142, 280.2292, 280.2024, 280.1755, 280.1487, 280.1218, 280.095, 
    280.0684, 280.0544, 280.0405, 280.0264, 280.0125, 279.9985, 279.9846, 
    279.9707, 279.9646, 279.9919, 280.0193, 280.0466, 280.074, 280.1013, 
    280.1265, 280.1348, 280.1431, 280.1514, 280.1597, 280.168, 280.1763, 
    280.1846, 280.1826, 280.1104, 280.0378, 279.9653, 279.8928, 279.8206, 
    279.7483, 279.6765, 279.6047, 279.533, 279.4612, 279.3894, 279.3176, 
    279.2458, 279.1748, 279.1179, 279.061, 279.0042, 278.9473, 278.8901, 
    278.8357, 278.7859, 278.7358, 278.686, 278.636, 278.5862, 278.5361, 
    278.4863, 278.4363, 278.4407, 278.4448, 278.4492, 278.4534, 278.4575, 
    278.4666, 278.481, 278.4954, 278.5098, 278.5242, 278.5386, 278.553, 
    278.5674, 278.582, 278.6299, 278.6799, 278.7302, 278.7803, 278.8306, 
    278.8743, 278.9133, 278.9524, 278.9917, 279.0308, 279.0698,
  276.5217, 276.5356, 276.5542, 276.5815, 276.6091, 276.6367, 276.6643, 
    276.6904, 276.707, 276.7236, 276.7402, 276.7568, 276.7734, 276.7903, 
    276.8069, 276.8235, 276.8445, 276.8706, 276.897, 276.9233, 276.9495, 
    276.979, 277.0552, 277.1316, 277.208, 277.2842, 277.3606, 277.437, 
    277.5134, 277.5896, 277.6638, 277.7366, 277.8091, 277.8818, 277.9543, 
    278.0271, 278.0723, 278.1174, 278.1626, 278.2078, 278.2529, 278.2981, 
    278.3433, 278.3884, 278.449, 278.5166, 278.5842, 278.6519, 278.7197, 
    278.7874, 278.8516, 278.9155, 278.9795, 279.0437, 279.1077, 279.1716, 
    279.2356, 279.2998, 279.3801, 279.4651, 279.5498, 279.6348, 279.7195, 
    279.8042, 279.9158, 280.0308, 280.146, 280.2612, 280.3762, 280.4915, 
    280.6067, 280.7217, 280.7651, 280.801, 280.8367, 280.8723, 280.9082, 
    280.9438, 280.9883, 281.0347, 281.0811, 281.1274, 281.1738, 281.2202, 
    281.2668, 281.3137, 281.4021, 281.4907, 281.5791, 281.6677, 281.7561, 
    281.8445, 281.8955, 281.9338, 281.9724, 282.0107, 282.0491, 282.0874, 
    282.126, 282.1606, 282.1709, 282.1809, 282.1909, 282.2009, 282.2109, 
    282.2212, 282.1582, 282.062, 281.9658, 281.8699, 281.7737, 281.6775, 
    281.5813, 281.4841, 281.3835, 281.283, 281.1821, 281.0815, 280.981, 
    280.8801, 280.8186, 280.7805, 280.7424, 280.7043, 280.6663, 280.6282, 
    280.5898, 280.5632, 280.5576, 280.552, 280.5464, 280.5408, 280.5352, 
    280.5293, 280.5579, 280.6125, 280.6675, 280.7224, 280.7771, 280.832, 
    280.887, 280.9412, 280.9949, 281.0486, 281.1023, 281.156, 281.2097, 
    281.2634, 281.3013, 281.3237, 281.3459, 281.3682, 281.3904, 281.4126, 
    281.4348, 281.447, 281.4517, 281.4563, 281.4609, 281.4658, 281.4705, 
    281.4751, 281.4873, 281.5095, 281.5315, 281.5535, 281.5754, 281.5977, 
    281.6196, 281.6375, 281.6533, 281.6692, 281.6851, 281.7009, 281.7168, 
    281.7327, 281.7422, 281.7415, 281.7407, 281.74, 281.7393, 281.7385, 
    281.7378, 281.728, 281.7161, 281.7041, 281.6921, 281.6802, 281.6682, 
    281.6562, 281.6155, 281.5112, 281.4072, 281.303, 281.199, 281.0947, 
    280.9907, 280.8962, 280.8027, 280.7092, 280.616, 280.5225, 280.429, 
    280.3357, 280.2583, 280.23, 280.2017, 280.1731, 280.1448, 280.1165, 
    280.0886, 280.0898, 280.0913, 280.0925, 280.0938, 280.0952, 280.0964, 
    280.0979, 280.1057, 280.1418, 280.1777, 280.2139, 280.2498, 280.2859, 
    280.3162, 280.3086, 280.3008, 280.293, 280.2852, 280.2773, 280.2698, 
    280.262, 280.2456, 280.1699, 280.0945, 280.0188, 279.9431, 279.8677, 
    279.7925, 279.7183, 279.6443, 279.5701, 279.4961, 279.4219, 279.3479, 
    279.2737, 279.2004, 279.1389, 279.0771, 279.0156, 278.9541, 278.8923, 
    278.8364, 278.791, 278.7454, 278.7, 278.6545, 278.6089, 278.5635, 
    278.5181, 278.4724, 278.4724, 278.4724, 278.4727, 278.4727, 278.4727, 
    278.4834, 278.5068, 278.5303, 278.5537, 278.5769, 278.6003, 278.6238, 
    278.6472, 278.6707, 278.7222, 278.7756, 278.8291, 278.8823, 278.9358, 
    278.9746, 279.0027, 279.0308, 279.0588, 279.0869, 279.115,
  276.4854, 276.4897, 276.5017, 276.5276, 276.5535, 276.5793, 276.6052, 
    276.6301, 276.6472, 276.6643, 276.6814, 276.6985, 276.7156, 276.7327, 
    276.7495, 276.7666, 276.7908, 276.8228, 276.855, 276.8872, 276.9192, 
    276.9541, 277.0266, 277.0994, 277.1721, 277.2449, 277.3176, 277.3901, 
    277.4629, 277.5356, 277.605, 277.6719, 277.7388, 277.8057, 277.8726, 
    277.9395, 277.9841, 278.0288, 278.0735, 278.1182, 278.1628, 278.2075, 
    278.2522, 278.2969, 278.3655, 278.4453, 278.5251, 278.605, 278.6848, 
    278.7646, 278.8416, 278.9185, 278.9954, 279.0723, 279.1492, 279.2261, 
    279.303, 279.3799, 279.4824, 279.5918, 279.7012, 279.8108, 279.9202, 
    280.0295, 280.1604, 280.2944, 280.4285, 280.5625, 280.6965, 280.8306, 
    280.9644, 281.0984, 281.1204, 281.1299, 281.1396, 281.1494, 281.1589, 
    281.1687, 281.1855, 281.2039, 281.2222, 281.2405, 281.2588, 281.2771, 
    281.2957, 281.3149, 281.3989, 281.4832, 281.5674, 281.6516, 281.7356, 
    281.8198, 281.8735, 281.9172, 281.9609, 282.0044, 282.0481, 282.0918, 
    282.1353, 282.1733, 282.1726, 282.1719, 282.1711, 282.1704, 282.1697, 
    282.1689, 282.1091, 282.0222, 281.9355, 281.8489, 281.7622, 281.6755, 
    281.5886, 281.5002, 281.4065, 281.3127, 281.2188, 281.125, 281.0312, 
    280.9375, 280.8752, 280.832, 280.7888, 280.7456, 280.7026, 280.6594, 
    280.6162, 280.5908, 280.5984, 280.6062, 280.6138, 280.6213, 280.6292, 
    280.6367, 280.6719, 280.7285, 280.7852, 280.8418, 280.8984, 280.9551, 
    281.0117, 281.0676, 281.1226, 281.1772, 281.2322, 281.2871, 281.3418, 
    281.3967, 281.439, 281.4683, 281.4976, 281.5271, 281.5564, 281.5857, 
    281.615, 281.6289, 281.6306, 281.6326, 281.6345, 281.6365, 281.6384, 
    281.6404, 281.6484, 281.6643, 281.6804, 281.6963, 281.7124, 281.7283, 
    281.7441, 281.7537, 281.76, 281.7664, 281.7727, 281.7791, 281.7852, 
    281.7915, 281.793, 281.7856, 281.7786, 281.7715, 281.7644, 281.7571, 
    281.75, 281.729, 281.7043, 281.6794, 281.6548, 281.6301, 281.6055, 
    281.5808, 281.5327, 281.4333, 281.334, 281.2346, 281.1353, 281.0359, 
    280.9368, 280.8525, 280.77, 280.6873, 280.6047, 280.5222, 280.4395, 
    280.3569, 280.2876, 280.2576, 280.2278, 280.1978, 280.1677, 280.1379, 
    280.1089, 280.1255, 280.1421, 280.1587, 280.1753, 280.1919, 280.2083, 
    280.2249, 280.2468, 280.2915, 280.3362, 280.3809, 280.4255, 280.4702, 
    280.5061, 280.4824, 280.4585, 280.4346, 280.4109, 280.387, 280.363, 
    280.3394, 280.3086, 280.2297, 280.1511, 280.0723, 279.9934, 279.9148, 
    279.8364, 279.7603, 279.6838, 279.6074, 279.531, 279.4546, 279.3782, 
    279.3018, 279.2261, 279.1597, 279.0935, 279.0271, 278.9609, 278.8945, 
    278.8372, 278.7961, 278.7551, 278.7139, 278.6729, 278.6318, 278.5908, 
    278.5498, 278.5085, 278.5044, 278.5002, 278.4961, 278.4917, 278.4875, 
    278.5002, 278.5327, 278.5649, 278.5974, 278.6299, 278.6621, 278.6946, 
    278.7268, 278.7593, 278.8145, 278.8711, 278.9277, 278.9846, 279.0413, 
    279.0752, 279.092, 279.1091, 279.126, 279.1431, 279.1602,
  276.449, 276.4441, 276.4492, 276.4734, 276.4978, 276.522, 276.5464, 
    276.5698, 276.5874, 276.6047, 276.6223, 276.6399, 276.6575, 276.6748, 
    276.6924, 276.71, 276.7368, 276.7749, 276.813, 276.8511, 276.8892, 
    276.929, 276.998, 277.0671, 277.1362, 277.2053, 277.2744, 277.3435, 
    277.4126, 277.4817, 277.5461, 277.6074, 277.6685, 277.7297, 277.7908, 
    277.8521, 277.8962, 277.9402, 277.9844, 278.0286, 278.0728, 278.1169, 
    278.1611, 278.2053, 278.282, 278.3738, 278.4658, 278.5579, 278.6499, 
    278.7419, 278.8318, 278.9214, 279.0112, 279.1011, 279.1907, 279.2805, 
    279.3701, 279.46, 279.5847, 279.7188, 279.8528, 279.9868, 280.1208, 
    280.2549, 280.4053, 280.5581, 280.7109, 280.8638, 281.0166, 281.1694, 
    281.3223, 281.4751, 281.4753, 281.459, 281.4426, 281.4263, 281.4099, 
    281.3936, 281.3826, 281.373, 281.3633, 281.3535, 281.3438, 281.3342, 
    281.3245, 281.3159, 281.3958, 281.4756, 281.5554, 281.6355, 281.7153, 
    281.7952, 281.8518, 281.9006, 281.9495, 281.9983, 282.0471, 282.0959, 
    282.1448, 282.186, 282.1743, 282.1628, 282.1514, 282.1399, 282.1282, 
    282.1167, 282.0601, 281.9827, 281.9053, 281.8281, 281.7507, 281.6733, 
    281.5959, 281.5164, 281.4294, 281.3425, 281.2556, 281.1685, 281.0815, 
    280.9946, 280.9319, 280.8835, 280.8354, 280.7871, 280.739, 280.6907, 
    280.6426, 280.6184, 280.6394, 280.6604, 280.6812, 280.7021, 280.7231, 
    280.7441, 280.7861, 280.8447, 280.9031, 280.9614, 281.0198, 281.0784, 
    281.1367, 281.1941, 281.25, 281.3062, 281.3621, 281.4182, 281.4741, 
    281.53, 281.5764, 281.6128, 281.6494, 281.686, 281.7224, 281.759, 
    281.7954, 281.8105, 281.8098, 281.8088, 281.8081, 281.8074, 281.8064, 
    281.8057, 281.8093, 281.8193, 281.8293, 281.8391, 281.8491, 281.8589, 
    281.8689, 281.8699, 281.8667, 281.8633, 281.8601, 281.8569, 281.8538, 
    281.8506, 281.8435, 281.8298, 281.8164, 281.803, 281.7893, 281.7759, 
    281.7625, 281.7297, 281.6924, 281.655, 281.6174, 281.5801, 281.5427, 
    281.5051, 281.45, 281.3555, 281.2607, 281.1663, 281.0718, 280.9773, 
    280.8828, 280.8088, 280.7371, 280.6653, 280.5935, 280.5217, 280.4502, 
    280.3784, 280.3167, 280.2852, 280.2537, 280.2224, 280.1909, 280.1594, 
    280.1292, 280.1609, 280.1929, 280.2246, 280.2566, 280.2883, 280.3203, 
    280.3521, 280.3879, 280.4414, 280.4946, 280.5481, 280.6013, 280.6548, 
    280.696, 280.656, 280.6162, 280.5764, 280.5364, 280.4966, 280.4565, 
    280.4167, 280.3716, 280.2896, 280.2078, 280.1257, 280.0437, 279.9619, 
    279.8806, 279.802, 279.7234, 279.6445, 279.5659, 279.4873, 279.4084, 
    279.3298, 279.2517, 279.1807, 279.1096, 279.0386, 278.9678, 278.8967, 
    278.8379, 278.8013, 278.7646, 278.728, 278.6914, 278.6548, 278.6179, 
    278.5813, 278.5447, 278.5364, 278.5278, 278.5195, 278.511, 278.5024, 
    278.5171, 278.5586, 278.5999, 278.6411, 278.6826, 278.7239, 278.7654, 
    278.8066, 278.8479, 278.9067, 278.9668, 279.0266, 279.0867, 279.1465, 
    279.1755, 279.1814, 279.1873, 279.1934, 279.1992, 279.2051,
  276.4126, 276.3982, 276.3967, 276.4194, 276.4421, 276.4648, 276.4873, 
    276.5095, 276.5273, 276.5454, 276.5635, 276.5813, 276.5994, 276.6172, 
    276.6353, 276.6533, 276.6831, 276.7271, 276.771, 276.8149, 276.8589, 
    276.9041, 276.9695, 277.0349, 277.1003, 277.1658, 277.2312, 277.2966, 
    277.3621, 277.4277, 277.4873, 277.5427, 277.5981, 277.6536, 277.709, 
    277.7644, 277.8081, 277.8518, 277.8953, 277.939, 277.9827, 278.0264, 
    278.0698, 278.1135, 278.1982, 278.3025, 278.4067, 278.5107, 278.615, 
    278.7192, 278.8218, 278.9243, 279.0271, 279.1296, 279.2322, 279.3347, 
    279.4375, 279.54, 279.687, 279.8457, 280.0042, 280.1628, 280.3215, 
    280.4802, 280.6501, 280.8218, 280.9934, 281.165, 281.3369, 281.5085, 
    281.6802, 281.8518, 281.8303, 281.7878, 281.7456, 281.7031, 281.6609, 
    281.6184, 281.5798, 281.542, 281.5044, 281.4666, 281.4287, 281.3911, 
    281.3533, 281.3171, 281.3926, 281.4683, 281.5437, 281.6194, 281.6948, 
    281.7703, 281.8298, 281.8838, 281.938, 281.9919, 282.0459, 282.1001, 
    282.1541, 282.1985, 282.1763, 282.1538, 282.1316, 282.1091, 282.0869, 
    282.0645, 282.011, 281.9429, 281.875, 281.8071, 281.7393, 281.6714, 
    281.6033, 281.5325, 281.4524, 281.3723, 281.2922, 281.2122, 281.1318, 
    281.0518, 280.9885, 280.9351, 280.8818, 280.8286, 280.7754, 280.7219, 
    280.6687, 280.646, 280.6802, 280.7146, 280.7488, 280.783, 280.8171, 
    280.8516, 280.9004, 280.9607, 281.0208, 281.0811, 281.1414, 281.2014, 
    281.2617, 281.3206, 281.3777, 281.4348, 281.4919, 281.5491, 281.6064, 
    281.6636, 281.7139, 281.7576, 281.8013, 281.845, 281.8884, 281.9321, 
    281.9758, 281.9924, 281.9888, 281.9854, 281.9817, 281.978, 281.9744, 
    281.9707, 281.9705, 281.9744, 281.9783, 281.9819, 281.9858, 281.9897, 
    281.9937, 281.9861, 281.9734, 281.9604, 281.9478, 281.9351, 281.9221, 
    281.9094, 281.894, 281.874, 281.8542, 281.8342, 281.8145, 281.7944, 
    281.7747, 281.7307, 281.6804, 281.6304, 281.5801, 281.53, 281.4797, 
    281.4297, 281.3672, 281.2773, 281.1877, 281.0979, 281.0083, 280.9185, 
    280.8289, 280.7651, 280.7043, 280.6433, 280.5825, 280.5215, 280.4607, 
    280.3997, 280.3457, 280.3127, 280.2798, 280.2468, 280.2139, 280.1809, 
    280.1494, 280.1965, 280.2437, 280.2908, 280.3379, 280.385, 280.4321, 
    280.4792, 280.5291, 280.5911, 280.6531, 280.7151, 280.7771, 280.8391, 
    280.886, 280.8298, 280.7739, 280.718, 280.6621, 280.606, 280.55, 
    280.4941, 280.4346, 280.3494, 280.2642, 280.1792, 280.094, 280.009, 
    279.9248, 279.8438, 279.7629, 279.6819, 279.6008, 279.5198, 279.4387, 
    279.3579, 279.2771, 279.2014, 279.126, 279.0503, 278.9746, 278.8989, 
    278.8386, 278.8064, 278.7742, 278.7419, 278.7097, 278.6775, 278.6453, 
    278.613, 278.5808, 278.5681, 278.5554, 278.543, 278.5303, 278.5176, 
    278.5339, 278.5845, 278.6348, 278.6851, 278.7354, 278.7856, 278.8359, 
    278.8862, 278.9368, 278.999, 279.0623, 279.1255, 279.1887, 279.252, 
    279.2759, 279.2708, 279.2656, 279.2605, 279.2554, 279.2502,
  276.3762, 276.3525, 276.3442, 276.3652, 276.3865, 276.4075, 276.4285, 
    276.4492, 276.4675, 276.4861, 276.5044, 276.5229, 276.5413, 276.5596, 
    276.5781, 276.5964, 276.6292, 276.6792, 276.729, 276.7788, 276.8286, 
    276.8792, 276.9409, 277.0027, 277.0647, 277.1265, 277.1882, 277.25, 
    277.3118, 277.3735, 277.4285, 277.4783, 277.5278, 277.5776, 277.6272, 
    277.677, 277.72, 277.7632, 277.8064, 277.8494, 277.8926, 277.9355, 
    277.9788, 278.022, 278.1147, 278.2312, 278.3474, 278.4639, 278.5801, 
    278.6965, 278.812, 278.9275, 279.0427, 279.1582, 279.2737, 279.3892, 
    279.5046, 279.6201, 279.7893, 279.9724, 280.1558, 280.3389, 280.5222, 
    280.7053, 280.895, 281.0854, 281.2759, 281.4666, 281.657, 281.8474, 
    282.0378, 282.2285, 282.1853, 282.1169, 282.0486, 281.9802, 281.9119, 
    281.8433, 281.7771, 281.7112, 281.6455, 281.5796, 281.5137, 281.448, 
    281.3821, 281.3181, 281.3894, 281.4607, 281.532, 281.603, 281.6743, 
    281.7456, 281.8079, 281.8672, 281.9263, 281.9856, 282.0449, 282.1042, 
    282.1633, 282.2112, 282.178, 282.1448, 282.1118, 282.0786, 282.0454, 
    282.0125, 281.9619, 281.9033, 281.8447, 281.7864, 281.7278, 281.6692, 
    281.6108, 281.5486, 281.4753, 281.4021, 281.3289, 281.2556, 281.1821, 
    281.1089, 281.0449, 280.9866, 280.9282, 280.8701, 280.8118, 280.7534, 
    280.6951, 280.6736, 280.7212, 280.7686, 280.8162, 280.8638, 280.9114, 
    280.959, 281.0146, 281.0767, 281.1387, 281.2007, 281.2627, 281.3247, 
    281.3867, 281.447, 281.5054, 281.5635, 281.6218, 281.6802, 281.7385, 
    281.7969, 281.8513, 281.9021, 281.9529, 282.0037, 282.0544, 282.1055, 
    282.1562, 282.1743, 282.168, 282.1616, 282.1553, 282.1487, 282.1423, 
    282.136, 282.1316, 282.1294, 282.127, 282.1248, 282.1226, 282.1204, 
    282.1182, 282.1023, 282.0798, 282.0576, 282.0354, 282.0129, 281.9907, 
    281.9685, 281.9446, 281.9182, 281.8921, 281.8657, 281.8394, 281.8132, 
    281.7869, 281.7314, 281.6687, 281.6057, 281.5427, 281.48, 281.417, 
    281.3542, 281.2844, 281.1995, 281.1145, 281.0295, 280.9446, 280.8599, 
    280.7749, 280.7214, 280.6714, 280.6213, 280.5713, 280.5212, 280.4712, 
    280.4211, 280.375, 280.3403, 280.3059, 280.2715, 280.2371, 280.2024, 
    280.1697, 280.2319, 280.2944, 280.3567, 280.4192, 280.4814, 280.5439, 
    280.6062, 280.6702, 280.741, 280.8115, 280.8823, 280.9529, 281.0234, 
    281.0759, 281.0037, 280.9316, 280.8596, 280.7876, 280.7156, 280.6436, 
    280.5715, 280.4973, 280.4092, 280.3208, 280.2327, 280.1443, 280.0562, 
    279.969, 279.8857, 279.8025, 279.719, 279.6357, 279.5525, 279.4692, 
    279.3857, 279.3027, 279.2224, 279.1421, 279.0618, 278.9814, 278.9011, 
    278.8394, 278.8115, 278.7837, 278.7559, 278.728, 278.7004, 278.6726, 
    278.6448, 278.6169, 278.6001, 278.5833, 278.5664, 278.5493, 278.5325, 
    278.551, 278.6101, 278.6694, 278.7288, 278.7881, 278.8474, 278.9067, 
    278.9661, 279.0254, 279.0913, 279.158, 279.2244, 279.2908, 279.3574, 
    279.3762, 279.3601, 279.344, 279.3276, 279.3115, 279.2954,
  276.3398, 276.3069, 276.292, 276.3113, 276.3306, 276.3501, 276.3694, 
    276.3889, 276.4077, 276.4265, 276.4453, 276.4644, 276.4832, 276.502, 
    276.521, 276.5398, 276.5754, 276.6311, 276.687, 276.7427, 276.7983, 
    276.8542, 276.9124, 276.9705, 277.0288, 277.0869, 277.145, 277.2034, 
    277.2615, 277.3196, 277.3696, 277.4136, 277.4575, 277.5015, 277.5454, 
    277.5894, 277.6321, 277.6746, 277.7173, 277.7598, 277.8025, 277.845, 
    277.8877, 277.9302, 278.0312, 278.1597, 278.2881, 278.4167, 278.5452, 
    278.6736, 278.802, 278.9304, 279.0586, 279.187, 279.3152, 279.4436, 
    279.572, 279.7002, 279.8914, 280.0994, 280.3071, 280.5149, 280.7229, 
    280.9307, 281.1399, 281.3491, 281.5586, 281.7678, 281.9771, 282.1865, 
    282.3958, 282.6052, 282.5403, 282.4458, 282.3516, 282.2571, 282.1626, 
    282.0684, 281.9744, 281.8804, 281.7866, 281.6926, 281.5986, 281.5049, 
    281.4109, 281.3193, 281.3862, 281.4531, 281.52, 281.5869, 281.6541, 
    281.7209, 281.7859, 281.8503, 281.9148, 281.9795, 282.0439, 282.1084, 
    282.1729, 282.2236, 282.1797, 282.1357, 282.092, 282.0481, 282.0042, 
    281.9602, 281.9126, 281.8635, 281.8145, 281.7654, 281.7163, 281.6672, 
    281.6182, 281.5649, 281.4983, 281.4319, 281.3655, 281.2991, 281.2327, 
    281.166, 281.1016, 281.0381, 280.9749, 280.9114, 280.8481, 280.7847, 
    280.7212, 280.7012, 280.762, 280.8228, 280.8838, 280.9446, 281.0054, 
    281.0662, 281.1287, 281.1926, 281.2563, 281.3201, 281.384, 281.4478, 
    281.5115, 281.5735, 281.6328, 281.6924, 281.7517, 281.8113, 281.8708, 
    281.9302, 281.989, 282.0469, 282.1047, 282.1626, 282.2207, 282.2786, 
    282.3364, 282.3562, 282.3469, 282.3379, 282.3286, 282.3196, 282.3105, 
    282.3013, 282.2925, 282.2842, 282.2759, 282.2676, 282.2595, 282.2512, 
    282.2429, 282.2185, 282.1865, 282.1548, 282.1228, 282.0911, 282.0591, 
    282.0273, 281.9951, 281.9624, 281.9299, 281.8972, 281.8645, 281.8318, 
    281.7991, 281.7324, 281.6567, 281.5811, 281.5056, 281.4299, 281.3542, 
    281.2786, 281.2017, 281.1216, 281.0413, 280.9612, 280.8811, 280.801, 
    280.7209, 280.6777, 280.6387, 280.5994, 280.5601, 280.521, 280.4817, 
    280.4426, 280.4041, 280.3682, 280.332, 280.2959, 280.26, 280.2239, 
    280.1899, 280.2676, 280.3452, 280.4229, 280.5005, 280.5781, 280.6558, 
    280.7334, 280.8113, 280.8906, 280.97, 281.0493, 281.1287, 281.208, 
    281.2656, 281.1775, 281.0896, 281.0015, 280.9133, 280.8252, 280.7371, 
    280.6489, 280.5603, 280.469, 280.3774, 280.2861, 280.1946, 280.1033, 
    280.0132, 279.9275, 279.842, 279.7563, 279.6707, 279.5852, 279.4995, 
    279.4138, 279.3284, 279.2434, 279.1582, 279.0732, 278.9883, 278.9033, 
    278.8401, 278.8167, 278.7932, 278.77, 278.7466, 278.7231, 278.7, 
    278.6765, 278.6531, 278.6321, 278.6108, 278.5898, 278.5686, 278.5474, 
    278.5679, 278.636, 278.7043, 278.7727, 278.8408, 278.9092, 278.9775, 
    279.0457, 279.114, 279.1836, 279.2534, 279.3232, 279.3931, 279.4626, 
    279.4768, 279.4495, 279.4221, 279.395, 279.3677, 279.3406,
  276.3293, 276.2959, 276.2803, 276.2983, 276.3164, 276.3345, 276.3525, 
    276.3706, 276.3887, 276.4067, 276.4248, 276.4429, 276.4607, 276.4788, 
    276.4968, 276.5149, 276.5532, 276.616, 276.6785, 276.741, 276.8037, 
    276.8662, 276.929, 276.9915, 277.054, 277.1167, 277.1792, 277.2417, 
    277.3044, 277.3669, 277.418, 277.4604, 277.5027, 277.5449, 277.5874, 
    277.6296, 277.6721, 277.7144, 277.7566, 277.7991, 277.8413, 277.8838, 
    277.926, 277.9683, 278.0691, 278.1973, 278.3252, 278.4534, 278.5815, 
    278.7097, 278.8379, 278.9661, 279.0942, 279.2222, 279.3503, 279.4785, 
    279.6067, 279.7349, 279.9326, 280.1489, 280.3652, 280.5815, 280.7979, 
    281.0139, 281.2302, 281.4465, 281.6628, 281.8792, 282.0955, 282.3118, 
    282.5278, 282.7441, 282.6829, 282.5916, 282.5002, 282.4089, 282.3176, 
    282.2263, 282.135, 282.0437, 281.9524, 281.8611, 281.7698, 281.6785, 
    281.5872, 281.4978, 281.5469, 281.5959, 281.6448, 281.6938, 281.7429, 
    281.7917, 281.8408, 281.8899, 281.9387, 281.9878, 282.0369, 282.0859, 
    282.1348, 282.1724, 282.1306, 282.0886, 282.0469, 282.0049, 281.9631, 
    281.9211, 281.8794, 281.8376, 281.7957, 281.7539, 281.7119, 281.6702, 
    281.6282, 281.582, 281.5225, 281.4629, 281.4031, 281.3435, 281.2839, 
    281.2241, 281.1646, 281.105, 281.0452, 280.9856, 280.926, 280.8662, 
    280.8066, 280.7898, 280.8533, 280.9165, 280.98, 281.0432, 281.1067, 
    281.1702, 281.2334, 281.2969, 281.3601, 281.4236, 281.4868, 281.5503, 
    281.6135, 281.6746, 281.7329, 281.791, 281.8494, 281.9077, 281.9658, 
    282.0242, 282.0825, 282.1406, 282.199, 282.2573, 282.3154, 282.3738, 
    282.4321, 282.4524, 282.4443, 282.4365, 282.4285, 282.4204, 282.4124, 
    282.4045, 282.3965, 282.3884, 282.3804, 282.3723, 282.3645, 282.3564, 
    282.3484, 282.3198, 282.2812, 282.2429, 282.2046, 282.1663, 282.1279, 
    282.0896, 282.0513, 282.0129, 281.9746, 281.9363, 281.8979, 281.8596, 
    281.8213, 281.7507, 281.6719, 281.593, 281.5139, 281.4351, 281.3562, 
    281.2773, 281.1985, 281.1194, 281.0405, 280.9617, 280.8828, 280.8037, 
    280.7249, 280.6877, 280.6548, 280.6218, 280.5889, 280.5559, 280.5229, 
    280.49, 280.457, 280.4241, 280.3911, 280.3582, 280.3252, 280.2922, 
    280.2612, 280.3342, 280.4075, 280.4805, 280.5537, 280.6267, 280.7, 
    280.7729, 280.8462, 280.9192, 280.9924, 281.0654, 281.1384, 281.2117, 
    281.2642, 281.1775, 281.0906, 281.0039, 280.9172, 280.8303, 280.7437, 
    280.6567, 280.5701, 280.4834, 280.3965, 280.3098, 280.2231, 280.1362, 
    280.05, 279.9658, 279.8813, 279.7971, 279.7126, 279.6282, 279.5439, 
    279.4595, 279.375, 279.2908, 279.2063, 279.1221, 279.0376, 278.9531, 
    278.8943, 278.8823, 278.8701, 278.8582, 278.8462, 278.834, 278.822, 
    278.8101, 278.7979, 278.7859, 278.7739, 278.7617, 278.7498, 278.7378, 
    278.7549, 278.8059, 278.8569, 278.908, 278.959, 279.01, 279.061, 
    279.1121, 279.1631, 279.2141, 279.2651, 279.3162, 279.3672, 279.4182, 
    279.4243, 279.3972, 279.3704, 279.3433, 279.3164, 279.2893,
  276.3279, 276.2971, 276.283, 276.2998, 276.3164, 276.3333, 276.3501, 
    276.3669, 276.3838, 276.4004, 276.4172, 276.4341, 276.4509, 276.4675, 
    276.4844, 276.5012, 276.5422, 276.6121, 276.6816, 276.7515, 276.8213, 
    276.8911, 276.9609, 277.0308, 277.1006, 277.1702, 277.24, 277.3098, 
    277.3796, 277.4495, 277.5034, 277.5457, 277.5879, 277.6299, 277.6721, 
    277.7144, 277.7563, 277.7986, 277.8408, 277.8828, 277.925, 277.9673, 
    278.0093, 278.0515, 278.1489, 278.2725, 278.3958, 278.5193, 278.6426, 
    278.7661, 278.8894, 279.0129, 279.1365, 279.2598, 279.3833, 279.5066, 
    279.6301, 279.7537, 279.9526, 280.1719, 280.3909, 280.6099, 280.8291, 
    281.0481, 281.2673, 281.4863, 281.7053, 281.9246, 282.1436, 282.3628, 
    282.5818, 282.8008, 282.7517, 282.6736, 282.5955, 282.5176, 282.4395, 
    282.3613, 282.2832, 282.2051, 282.127, 282.0488, 281.9707, 281.8926, 
    281.8145, 281.7378, 281.7642, 281.7905, 281.8169, 281.8433, 281.8696, 
    281.896, 281.9224, 281.9487, 281.9751, 282.0015, 282.0278, 282.0542, 
    282.0803, 282.0991, 282.0637, 282.0283, 281.9929, 281.9575, 281.9224, 
    281.887, 281.8516, 281.8162, 281.7808, 281.7454, 281.7102, 281.6748, 
    281.6394, 281.5999, 281.5471, 281.4941, 281.4412, 281.3884, 281.3354, 
    281.2827, 281.2297, 281.177, 281.124, 281.0713, 281.0183, 280.9653, 
    280.9126, 280.8997, 280.9619, 281.0242, 281.0862, 281.1484, 281.2104, 
    281.2727, 281.3347, 281.397, 281.459, 281.5212, 281.5833, 281.6455, 
    281.7075, 281.7671, 281.8232, 281.8796, 281.9358, 281.9919, 282.0483, 
    282.1045, 282.1606, 282.217, 282.2732, 282.3296, 282.3857, 282.4419, 
    282.4983, 282.5193, 282.5137, 282.5081, 282.5027, 282.4971, 282.4915, 
    282.4861, 282.4805, 282.4751, 282.4695, 282.4639, 282.4585, 282.4529, 
    282.4475, 282.4158, 282.3721, 282.3281, 282.2844, 282.2407, 282.197, 
    282.1531, 282.1094, 282.0657, 282.022, 281.978, 281.9343, 281.8906, 
    281.8469, 281.7751, 281.6963, 281.6172, 281.5383, 281.4595, 281.3806, 
    281.3015, 281.2227, 281.1438, 281.0647, 280.9858, 280.907, 280.8281, 
    280.749, 280.7161, 280.6877, 280.6594, 280.6313, 280.603, 280.5747, 
    280.5464, 280.5183, 280.49, 280.4617, 280.4333, 280.4053, 280.377, 
    280.3501, 280.4119, 280.4736, 280.5354, 280.5972, 280.6589, 280.7205, 
    280.7822, 280.844, 280.9058, 280.9675, 281.0293, 281.0908, 281.1526, 
    281.1963, 281.1169, 281.0376, 280.958, 280.8787, 280.7993, 280.72, 
    280.6406, 280.5613, 280.4819, 280.4026, 280.3232, 280.2439, 280.1646, 
    280.0847, 280.0027, 279.9209, 279.8389, 279.7571, 279.675, 279.593, 
    279.5112, 279.4292, 279.3474, 279.2654, 279.1836, 279.1016, 279.0198, 
    278.9673, 278.969, 278.9705, 278.9722, 278.9739, 278.9756, 278.9773, 
    278.9788, 278.9805, 278.9822, 278.9839, 278.9856, 278.9871, 278.9888, 
    279.0012, 279.0259, 279.0505, 279.0752, 279.0996, 279.1243, 279.1489, 
    279.1736, 279.1982, 279.2229, 279.2476, 279.2722, 279.2969, 279.3215, 
    279.3188, 279.2961, 279.2734, 279.2505, 279.2278, 279.2051,
  276.3264, 276.2986, 276.2856, 276.301, 276.3167, 276.332, 276.3477, 
    276.3633, 276.3787, 276.3943, 276.4097, 276.4253, 276.4409, 276.4563, 
    276.4719, 276.4873, 276.531, 276.6079, 276.6851, 276.762, 276.8389, 
    276.916, 276.9929, 277.0698, 277.147, 277.2239, 277.301, 277.3779, 
    277.4548, 277.532, 277.5889, 277.6309, 277.6729, 277.7148, 277.7568, 
    277.7988, 277.8408, 277.8828, 277.9248, 277.9668, 278.0088, 278.0508, 
    278.0928, 278.1348, 278.2288, 278.3477, 278.4663, 278.585, 278.7039, 
    278.8225, 278.9412, 279.0601, 279.1787, 279.2974, 279.4163, 279.5349, 
    279.6536, 279.7725, 279.9727, 280.1946, 280.4165, 280.6384, 280.8604, 
    281.0823, 281.3042, 281.5261, 281.748, 281.97, 282.1919, 282.4138, 
    282.6357, 282.8577, 282.8206, 282.7559, 282.6909, 282.626, 282.561, 
    282.4961, 282.4314, 282.3665, 282.3015, 282.2366, 282.1716, 282.1067, 
    282.042, 281.978, 281.9817, 281.9854, 281.989, 281.9927, 281.9963, 
    282.0002, 282.0039, 282.0076, 282.0112, 282.0149, 282.0186, 282.0225, 
    282.0261, 282.0256, 281.9968, 281.968, 281.9392, 281.9102, 281.8813, 
    281.8525, 281.8237, 281.7949, 281.7659, 281.7371, 281.7083, 281.6794, 
    281.6506, 281.6177, 281.5715, 281.5254, 281.4792, 281.4333, 281.3872, 
    281.3411, 281.2949, 281.2488, 281.2029, 281.1567, 281.1106, 281.0645, 
    281.0186, 281.0098, 281.0706, 281.1316, 281.1924, 281.2534, 281.3142, 
    281.3752, 281.436, 281.4971, 281.5579, 281.6189, 281.6797, 281.7407, 
    281.8015, 281.8594, 281.9136, 281.968, 282.0222, 282.0764, 282.1306, 
    282.1848, 282.239, 282.2932, 282.3474, 282.4016, 282.4561, 282.5103, 
    282.5645, 282.5859, 282.5828, 282.5798, 282.5767, 282.5737, 282.5708, 
    282.5676, 282.5647, 282.5615, 282.5586, 282.5554, 282.5525, 282.5493, 
    282.5464, 282.5117, 282.4626, 282.4136, 282.3643, 282.3152, 282.2659, 
    282.2168, 282.1675, 282.1184, 282.0691, 282.02, 281.9707, 281.9216, 
    281.8723, 281.7996, 281.7207, 281.6416, 281.5627, 281.4839, 281.4048, 
    281.3259, 281.2471, 281.168, 281.0891, 281.01, 280.9312, 280.8523, 
    280.7732, 280.7444, 280.7209, 280.6973, 280.6738, 280.6501, 280.6265, 
    280.603, 280.5793, 280.5559, 280.5322, 280.5085, 280.4851, 280.4614, 
    280.4392, 280.4895, 280.5398, 280.5903, 280.6406, 280.6909, 280.7412, 
    280.7915, 280.842, 280.8923, 280.9426, 280.9929, 281.0432, 281.0938, 
    281.1282, 281.0564, 280.9844, 280.9124, 280.8403, 280.7686, 280.6965, 
    280.6245, 280.5527, 280.4807, 280.4087, 280.3367, 280.2649, 280.1929, 
    280.1191, 280.0396, 279.9602, 279.8809, 279.8013, 279.7219, 279.6423, 
    279.563, 279.4834, 279.4041, 279.3245, 279.2451, 279.1658, 279.0862, 
    279.04, 279.0554, 279.0708, 279.0862, 279.1016, 279.1169, 279.1323, 
    279.1477, 279.1631, 279.1785, 279.1938, 279.2092, 279.2246, 279.24, 
    279.2473, 279.2456, 279.2439, 279.2422, 279.2405, 279.2388, 279.2371, 
    279.2354, 279.2336, 279.2319, 279.23, 279.2283, 279.2266, 279.2249, 
    279.2134, 279.1948, 279.1763, 279.1577, 279.1392, 279.1206,
  276.325, 276.2998, 276.2881, 276.3025, 276.3167, 276.3311, 276.3452, 
    276.3596, 276.3738, 276.3879, 276.4023, 276.4165, 276.4309, 276.4451, 
    276.4595, 276.4736, 276.5198, 276.604, 276.6882, 276.7725, 276.8567, 
    276.9409, 277.0249, 277.1091, 277.1934, 277.2776, 277.3618, 277.446, 
    277.5303, 277.6143, 277.6746, 277.7163, 277.7581, 277.7998, 277.8416, 
    277.8835, 277.9253, 277.967, 278.0088, 278.0505, 278.0925, 278.1343, 
    278.176, 278.2178, 278.3086, 278.4229, 278.5369, 278.6509, 278.7649, 
    278.8789, 278.9929, 279.1069, 279.2209, 279.335, 279.449, 279.563, 
    279.677, 279.791, 279.9927, 280.2175, 280.4421, 280.667, 280.8916, 
    281.1165, 281.3411, 281.5659, 281.7905, 282.0154, 282.24, 282.4648, 
    282.6895, 282.9143, 282.8896, 282.8379, 282.7861, 282.7344, 282.6829, 
    282.6311, 282.5793, 282.5276, 282.4761, 282.4243, 282.3726, 282.321, 
    282.2693, 282.218, 282.199, 282.1802, 282.1611, 282.1423, 282.1233, 
    282.1042, 282.0854, 282.0664, 282.0474, 282.0286, 282.0095, 281.9907, 
    281.9717, 281.9524, 281.9299, 281.9075, 281.8853, 281.8628, 281.8406, 
    281.8181, 281.7959, 281.7734, 281.7512, 281.7288, 281.7063, 281.6841, 
    281.6616, 281.6353, 281.5959, 281.5566, 281.5173, 281.478, 281.4387, 
    281.3994, 281.3601, 281.3208, 281.2815, 281.2422, 281.2029, 281.1636, 
    281.1243, 281.1196, 281.1792, 281.239, 281.2986, 281.3584, 281.418, 
    281.4778, 281.5374, 281.5972, 281.657, 281.7166, 281.7764, 281.8359, 
    281.8958, 281.9519, 282.0042, 282.0564, 282.1086, 282.1606, 282.2129, 
    282.2651, 282.3174, 282.3696, 282.4216, 282.4739, 282.5261, 282.5784, 
    282.6306, 282.6526, 282.6521, 282.6516, 282.6509, 282.6504, 282.6499, 
    282.6492, 282.6487, 282.6482, 282.6477, 282.647, 282.6465, 282.646, 
    282.6453, 282.6079, 282.5532, 282.4988, 282.4441, 282.3894, 282.335, 
    282.2803, 282.2256, 282.1711, 282.1165, 282.0618, 282.0073, 281.9526, 
    281.8979, 281.824, 281.7451, 281.666, 281.5872, 281.5081, 281.4292, 
    281.3503, 281.2712, 281.1924, 281.1133, 281.0344, 280.9553, 280.8765, 
    280.7974, 280.7729, 280.7539, 280.7351, 280.7163, 280.6973, 280.6785, 
    280.6594, 280.6406, 280.6218, 280.6028, 280.584, 280.5649, 280.5461, 
    280.5283, 280.5671, 280.6062, 280.645, 280.6841, 280.7229, 280.762, 
    280.801, 280.8398, 280.8789, 280.9177, 280.9568, 280.9956, 281.0347, 
    281.0603, 280.9956, 280.9312, 280.8667, 280.802, 280.7375, 280.6731, 
    280.6084, 280.5439, 280.4792, 280.4148, 280.3503, 280.2856, 280.2212, 
    280.1536, 280.0767, 279.9995, 279.9226, 279.8457, 279.7686, 279.6917, 
    279.6147, 279.5376, 279.4607, 279.3838, 279.3066, 279.2297, 279.1526, 
    279.113, 279.1421, 279.1711, 279.2002, 279.2292, 279.2583, 279.2874, 
    279.3167, 279.3457, 279.3748, 279.4038, 279.4329, 279.4619, 279.491, 
    279.4937, 279.4656, 279.4373, 279.4092, 279.3811, 279.353, 279.325, 
    279.2969, 279.2688, 279.2407, 279.2126, 279.1846, 279.1565, 279.1282, 
    279.1082, 279.0938, 279.0793, 279.0649, 279.0505, 279.0361,
  276.3235, 276.301, 276.2908, 276.3037, 276.3169, 276.3298, 276.3428, 
    276.356, 276.3689, 276.3818, 276.3948, 276.408, 276.4209, 276.4338, 
    276.4468, 276.46, 276.5088, 276.6001, 276.6914, 276.783, 276.8743, 
    276.9656, 277.0571, 277.1484, 277.2397, 277.3313, 277.4226, 277.5142, 
    277.6055, 277.6968, 277.76, 277.8015, 277.8433, 277.8848, 277.9265, 
    277.968, 278.0098, 278.0513, 278.0928, 278.1345, 278.176, 278.2178, 
    278.2593, 278.301, 278.3887, 278.4978, 278.6072, 278.7166, 278.8259, 
    278.9353, 279.0447, 279.1538, 279.2632, 279.3726, 279.4819, 279.5913, 
    279.7004, 279.8098, 280.0127, 280.2402, 280.4678, 280.6953, 280.9229, 
    281.1504, 281.3782, 281.6057, 281.8333, 282.0608, 282.2883, 282.5159, 
    282.7434, 282.9709, 282.9585, 282.9199, 282.8813, 282.843, 282.8044, 
    282.7661, 282.7275, 282.689, 282.6506, 282.6121, 282.5735, 282.5352, 
    282.4966, 282.458, 282.4165, 282.3748, 282.3333, 282.2917, 282.25, 
    282.2085, 282.1667, 282.1252, 282.0837, 282.042, 282.0005, 281.959, 
    281.9172, 281.8789, 281.863, 281.8472, 281.8313, 281.8154, 281.7996, 
    281.7837, 281.7681, 281.7522, 281.7363, 281.7205, 281.7046, 281.6887, 
    281.6729, 281.6531, 281.6206, 281.5879, 281.5554, 281.5229, 281.4905, 
    281.458, 281.4253, 281.3928, 281.3604, 281.3279, 281.2954, 281.2627, 
    281.2302, 281.2295, 281.2878, 281.3464, 281.4048, 281.4634, 281.522, 
    281.5803, 281.6389, 281.6973, 281.7559, 281.8142, 281.8728, 281.9312, 
    281.9897, 282.0444, 282.0945, 282.1448, 282.1948, 282.2451, 282.2952, 
    282.3455, 282.3958, 282.4458, 282.4961, 282.5461, 282.5964, 282.6465, 
    282.6968, 282.7192, 282.7212, 282.7231, 282.7251, 282.7271, 282.729, 
    282.731, 282.7329, 282.7346, 282.7366, 282.7385, 282.7405, 282.7424, 
    282.7444, 282.7039, 282.6438, 282.584, 282.5239, 282.4639, 282.4038, 
    282.3438, 282.2837, 282.2236, 282.1636, 282.1038, 282.0437, 281.9836, 
    281.9236, 281.8484, 281.7695, 281.6904, 281.6116, 281.5325, 281.4536, 
    281.3745, 281.2957, 281.2166, 281.1377, 281.0586, 280.9795, 280.9006, 
    280.8215, 280.8013, 280.7871, 280.7729, 280.7588, 280.7444, 280.7302, 
    280.7161, 280.7019, 280.6875, 280.6733, 280.6592, 280.645, 280.6306, 
    280.6172, 280.6448, 280.6724, 280.7, 280.7275, 280.7551, 280.7827, 
    280.8103, 280.8379, 280.8655, 280.8928, 280.9204, 280.948, 280.9756, 
    280.9922, 280.9351, 280.8779, 280.8208, 280.7637, 280.7065, 280.6494, 
    280.5923, 280.5352, 280.478, 280.4209, 280.3638, 280.3066, 280.2495, 
    280.1882, 280.1135, 280.0391, 279.9646, 279.8899, 279.8154, 279.741, 
    279.6663, 279.5918, 279.5173, 279.4429, 279.3682, 279.2937, 279.2192, 
    279.186, 279.2288, 279.2715, 279.3142, 279.3569, 279.3999, 279.4426, 
    279.4854, 279.5281, 279.571, 279.6138, 279.6565, 279.6992, 279.7422, 
    279.7397, 279.6853, 279.6309, 279.5764, 279.522, 279.4675, 279.4128, 
    279.3584, 279.304, 279.2495, 279.1951, 279.1406, 279.0862, 279.0317, 
    279.0027, 278.9924, 278.9824, 278.9722, 278.9619, 278.9519,
  276.322, 276.3022, 276.2935, 276.3052, 276.3169, 276.3286, 276.3403, 
    276.3521, 276.364, 276.3757, 276.3875, 276.3992, 276.4109, 276.4226, 
    276.4343, 276.446, 276.4976, 276.5962, 276.6948, 276.7932, 276.8918, 
    276.9905, 277.0891, 277.1877, 277.2864, 277.385, 277.4834, 277.582, 
    277.6807, 277.7793, 277.8455, 277.887, 277.9282, 277.9697, 278.0112, 
    278.0527, 278.094, 278.1355, 278.177, 278.2183, 278.2598, 278.3013, 
    278.3428, 278.384, 278.4685, 278.573, 278.6777, 278.7825, 278.887, 
    278.9917, 279.0962, 279.2009, 279.3054, 279.4102, 279.5146, 279.6194, 
    279.7241, 279.8286, 280.0327, 280.2632, 280.4934, 280.7239, 280.9543, 
    281.1846, 281.415, 281.6455, 281.8757, 282.1062, 282.3364, 282.5669, 
    282.7974, 283.0276, 283.0273, 283.002, 282.9768, 282.9514, 282.9263, 
    282.9009, 282.8757, 282.8503, 282.8252, 282.7998, 282.7744, 282.7493, 
    282.7239, 282.6982, 282.6338, 282.5696, 282.5054, 282.4412, 282.377, 
    282.3127, 282.2483, 282.1841, 282.1199, 282.0557, 281.9915, 281.9272, 
    281.8628, 281.8054, 281.7961, 281.7869, 281.7776, 281.7681, 281.7588, 
    281.7495, 281.74, 281.7307, 281.7214, 281.7122, 281.7026, 281.6934, 
    281.6841, 281.6707, 281.645, 281.6194, 281.5935, 281.5679, 281.542, 
    281.5164, 281.4907, 281.4648, 281.4392, 281.4133, 281.3877, 281.3618, 
    281.3362, 281.3394, 281.3967, 281.4539, 281.5112, 281.5684, 281.6257, 
    281.6829, 281.7402, 281.7974, 281.8547, 281.9119, 281.9692, 282.0264, 
    282.0837, 282.1367, 282.1851, 282.2332, 282.2812, 282.3293, 282.3777, 
    282.4258, 282.4739, 282.522, 282.5703, 282.6184, 282.6665, 282.7148, 
    282.7629, 282.7861, 282.7905, 282.7949, 282.7993, 282.8037, 282.8081, 
    282.8125, 282.8169, 282.8213, 282.8257, 282.8301, 282.8345, 282.8389, 
    282.8433, 282.8, 282.7346, 282.6692, 282.6038, 282.5381, 282.4727, 
    282.4072, 282.3418, 282.2764, 282.2109, 282.1455, 282.0801, 282.0146, 
    281.9492, 281.8728, 281.7939, 281.7148, 281.636, 281.5569, 281.4778, 
    281.3989, 281.3198, 281.241, 281.1619, 281.0828, 281.0039, 280.9248, 
    280.8457, 280.8298, 280.8203, 280.8108, 280.801, 280.7915, 280.782, 
    280.7725, 280.7629, 280.7534, 280.7439, 280.7344, 280.7249, 280.7153, 
    280.7063, 280.7224, 280.7385, 280.7549, 280.771, 280.7871, 280.8032, 
    280.8196, 280.8357, 280.8518, 280.8682, 280.8843, 280.9004, 280.9167, 
    280.9243, 280.8745, 280.825, 280.7751, 280.7253, 280.6755, 280.626, 
    280.5762, 280.5264, 280.4766, 280.427, 280.3772, 280.3274, 280.2778, 
    280.2227, 280.1506, 280.0784, 280.0063, 279.9343, 279.8623, 279.7903, 
    279.718, 279.646, 279.574, 279.502, 279.4297, 279.3577, 279.2856, 
    279.2588, 279.3154, 279.3718, 279.4282, 279.4849, 279.5413, 279.5977, 
    279.6543, 279.7107, 279.7671, 279.8237, 279.8801, 279.9368, 279.9932, 
    279.9861, 279.905, 279.8242, 279.7434, 279.6626, 279.5818, 279.501, 
    279.4202, 279.3394, 279.2585, 279.1775, 279.0967, 279.0159, 278.9351, 
    278.8972, 278.8914, 278.8853, 278.8794, 278.8735, 278.8674,
  276.3206, 276.3035, 276.2961, 276.3066, 276.3171, 276.3274, 276.3379, 
    276.3484, 276.3589, 276.3694, 276.3799, 276.3904, 276.4009, 276.4114, 
    276.4219, 276.4324, 276.4863, 276.5923, 276.698, 276.8037, 276.9097, 
    277.0154, 277.1211, 277.2271, 277.3328, 277.4385, 277.5444, 277.6501, 
    277.7561, 277.8618, 277.9309, 277.9722, 278.0134, 278.0547, 278.0959, 
    278.1372, 278.1785, 278.2197, 278.261, 278.3022, 278.3435, 278.3848, 
    278.426, 278.4673, 278.5483, 278.6482, 278.7483, 278.8481, 278.948, 
    279.0481, 279.1479, 279.2478, 279.3479, 279.4478, 279.5476, 279.6475, 
    279.7476, 279.8474, 280.0527, 280.2859, 280.519, 280.7524, 280.9856, 
    281.2188, 281.4519, 281.6851, 281.9185, 282.1516, 282.3848, 282.6179, 
    282.8511, 283.0845, 283.0962, 283.0842, 283.072, 283.0601, 283.0479, 
    283.0359, 283.0237, 283.0117, 282.9995, 282.9875, 282.9753, 282.9634, 
    282.9514, 282.9382, 282.8513, 282.7644, 282.6775, 282.5906, 282.5037, 
    282.4167, 282.3298, 282.2429, 282.156, 282.0691, 281.9822, 281.8955, 
    281.8086, 281.7322, 281.7292, 281.7266, 281.7236, 281.7207, 281.718, 
    281.7151, 281.7122, 281.7095, 281.7065, 281.7036, 281.7009, 281.698, 
    281.6951, 281.6885, 281.6694, 281.6506, 281.6316, 281.6128, 281.5938, 
    281.5747, 281.5559, 281.5369, 281.5178, 281.499, 281.48, 281.4609, 
    281.4421, 281.4492, 281.5054, 281.5613, 281.6174, 281.6733, 281.7295, 
    281.7854, 281.8416, 281.8975, 281.9536, 282.0095, 282.0657, 282.1218, 
    282.1777, 282.2292, 282.2754, 282.3215, 282.3677, 282.4138, 282.46, 
    282.5061, 282.5522, 282.5984, 282.6445, 282.6907, 282.7368, 282.783, 
    282.8291, 282.8528, 282.8596, 282.8665, 282.8735, 282.8804, 282.8872, 
    282.894, 282.9009, 282.908, 282.9148, 282.9216, 282.9285, 282.9353, 
    282.9424, 282.896, 282.8252, 282.7544, 282.6833, 282.6125, 282.5417, 
    282.4707, 282.3999, 282.3291, 282.2583, 282.1873, 282.1165, 282.0457, 
    281.9746, 281.8975, 281.8184, 281.7393, 281.6602, 281.5813, 281.5022, 
    281.4231, 281.3442, 281.2651, 281.186, 281.1072, 281.0281, 280.949, 
    280.8699, 280.8582, 280.8533, 280.8484, 280.8435, 280.8386, 280.834, 
    280.8291, 280.8242, 280.8193, 280.8145, 280.8096, 280.8047, 280.7998, 
    280.7952, 280.8, 280.8049, 280.8096, 280.8145, 280.8193, 280.824, 
    280.8289, 280.8337, 280.8384, 280.8433, 280.8481, 280.8528, 280.8577, 
    280.8564, 280.814, 280.7717, 280.7292, 280.687, 280.6448, 280.6023, 
    280.5601, 280.5176, 280.4753, 280.4331, 280.3906, 280.3484, 280.3059, 
    280.2571, 280.1875, 280.1179, 280.0483, 279.9788, 279.9089, 279.8394, 
    279.7698, 279.7002, 279.6306, 279.561, 279.4915, 279.4219, 279.3521, 
    279.3318, 279.4019, 279.4722, 279.5422, 279.6125, 279.6826, 279.7529, 
    279.823, 279.8933, 279.9634, 280.0337, 280.1038, 280.1741, 280.2441, 
    280.2322, 280.125, 280.0178, 279.9106, 279.8035, 279.696, 279.5889, 
    279.4817, 279.3745, 279.2673, 279.1602, 279.053, 278.9456, 278.8384, 
    278.792, 278.79, 278.7883, 278.7866, 278.7849, 278.783,
  276.354, 276.3423, 276.3384, 276.3501, 276.3618, 276.3735, 276.3853, 
    276.397, 276.4087, 276.4204, 276.4321, 276.4438, 276.4575, 276.4749, 
    276.4924, 276.5098, 276.5674, 276.6726, 276.7778, 276.8831, 276.9883, 
    277.0935, 277.1987, 277.304, 277.4092, 277.5144, 277.6194, 277.7246, 
    277.8296, 277.9348, 278.0059, 278.051, 278.0964, 278.1416, 278.1868, 
    278.2319, 278.2773, 278.3225, 278.3677, 278.4124, 278.457, 278.5015, 
    278.5459, 278.5903, 278.6699, 278.7659, 278.8621, 278.958, 279.0542, 
    279.1501, 279.2461, 279.3423, 279.4404, 279.5425, 279.6445, 279.7466, 
    279.8486, 279.9507, 280.1492, 280.3728, 280.5967, 280.8203, 281.0442, 
    281.2678, 281.4917, 281.7156, 281.9402, 282.165, 282.3899, 282.6147, 
    282.8396, 283.0645, 283.0928, 283.0999, 283.1072, 283.1143, 283.1213, 
    283.1287, 283.1357, 283.1238, 283.1028, 283.0818, 283.0608, 283.0398, 
    283.0186, 282.9966, 282.8992, 282.8018, 282.7043, 282.6067, 282.5093, 
    282.4119, 282.3188, 282.2344, 282.1497, 282.0652, 281.9807, 281.896, 
    281.8115, 281.7373, 281.7356, 281.7341, 281.7327, 281.731, 281.7295, 
    281.7278, 281.7236, 281.7197, 281.7156, 281.7114, 281.7073, 281.7031, 
    281.6992, 281.6917, 281.6731, 281.6545, 281.6362, 281.6177, 281.5991, 
    281.5867, 281.5771, 281.5676, 281.5581, 281.5486, 281.5391, 281.5295, 
    281.52, 281.5332, 281.5889, 281.6448, 281.7004, 281.7563, 281.8123, 
    281.8684, 281.9246, 281.9807, 282.0371, 282.0933, 282.1494, 282.2056, 
    282.2617, 282.314, 282.3608, 282.408, 282.4551, 282.5022, 282.5454, 
    282.5886, 282.6316, 282.6748, 282.718, 282.7612, 282.8042, 282.8474, 
    282.8906, 282.9143, 282.9233, 282.9324, 282.9414, 282.9438, 282.9436, 
    282.9431, 282.9426, 282.9421, 282.9417, 282.9412, 282.9407, 282.9404, 
    282.9399, 282.8904, 282.8179, 282.7456, 282.6743, 282.6052, 282.5359, 
    282.4666, 282.3975, 282.3281, 282.259, 282.1897, 282.1206, 282.0513, 
    281.9819, 281.908, 281.833, 281.7578, 281.6833, 281.6089, 281.5344, 
    281.46, 281.3855, 281.3108, 281.2363, 281.1619, 281.0874, 281.0129, 
    280.9385, 280.9255, 280.9189, 280.9126, 280.9062, 280.8999, 280.8936, 
    280.8872, 280.8809, 280.8745, 280.8684, 280.8621, 280.8557, 280.8494, 
    280.8433, 280.8413, 280.842, 280.8474, 280.8525, 280.8579, 280.8633, 
    280.8684, 280.8738, 280.8789, 280.8843, 280.8896, 280.8948, 280.9001, 
    280.9006, 280.8679, 280.8213, 280.7744, 280.7275, 280.6807, 280.634, 
    280.5872, 280.5403, 280.4934, 280.4468, 280.3999, 280.353, 280.3062, 
    280.2532, 280.1841, 280.1167, 280.0493, 279.9817, 279.9143, 279.8469, 
    279.7795, 279.7119, 279.6445, 279.5771, 279.5098, 279.4421, 279.3748, 
    279.3569, 279.4307, 279.5042, 279.5779, 279.6514, 279.7251, 279.7986, 
    279.8723, 279.946, 280.0195, 280.0933, 280.1667, 280.2405, 280.3137, 
    280.2878, 280.1707, 280.0537, 279.9368, 279.8198, 279.7029, 279.5857, 
    279.4688, 279.3518, 279.2349, 279.1177, 279.0007, 278.8838, 278.7759, 
    278.731, 278.7297, 278.7283, 278.7271, 278.7258, 278.7246,
  276.4016, 276.3958, 276.3967, 276.4106, 276.4246, 276.4385, 276.4524, 
    276.4663, 276.4805, 276.4944, 276.5083, 276.5222, 276.5408, 276.5684, 
    276.5962, 276.6238, 276.6851, 276.7866, 276.8882, 276.9897, 277.0913, 
    277.1926, 277.2942, 277.3958, 277.4973, 277.5989, 277.7002, 277.8013, 
    277.9026, 278.0039, 278.0767, 278.1274, 278.1782, 278.2292, 278.28, 
    278.3311, 278.3818, 278.4326, 278.4836, 278.5332, 278.5823, 278.6313, 
    278.6804, 278.7295, 278.8081, 278.9006, 278.9932, 279.0857, 279.178, 
    279.2705, 279.363, 279.4556, 279.553, 279.6599, 279.7671, 279.874, 
    279.981, 280.0881, 280.2761, 280.4854, 280.6948, 280.9043, 281.1138, 
    281.3232, 281.5325, 281.7419, 281.9539, 282.166, 282.3779, 282.5898, 
    282.802, 283.0139, 283.0605, 283.0894, 283.1182, 283.1467, 283.1755, 
    283.2043, 283.2332, 283.2161, 283.1772, 283.1384, 283.0996, 283.0608, 
    283.022, 282.9822, 282.8792, 282.7759, 282.6729, 282.5696, 282.4666, 
    282.3633, 282.2708, 282.1987, 282.1265, 282.0542, 281.9819, 281.9097, 
    281.8374, 281.7739, 281.7715, 281.769, 281.7668, 281.7644, 281.762, 
    281.7595, 281.751, 281.7427, 281.7341, 281.7256, 281.7173, 281.7087, 
    281.7002, 281.689, 281.6685, 281.6477, 281.6272, 281.6067, 281.5859, 
    281.5801, 281.5811, 281.5818, 281.5828, 281.5837, 281.5847, 281.5857, 
    281.5864, 281.6067, 281.6626, 281.7185, 281.7742, 281.8301, 281.8865, 
    281.9434, 282.0002, 282.0571, 282.1143, 282.1711, 282.228, 282.2849, 
    282.3418, 282.3953, 282.4446, 282.4939, 282.5432, 282.5923, 282.6321, 
    282.6719, 282.7117, 282.7515, 282.7913, 282.8311, 282.8706, 282.9104, 
    282.9502, 282.9736, 282.9846, 282.9958, 283.0068, 283.0024, 282.9907, 
    282.979, 282.9673, 282.9556, 282.9438, 282.9321, 282.9204, 282.9084, 
    282.8967, 282.8438, 282.7715, 282.6992, 282.6296, 282.5649, 282.5002, 
    282.4353, 282.3706, 282.3059, 282.2412, 282.1763, 282.1116, 282.0469, 
    281.9819, 281.9133, 281.8435, 281.7739, 281.7058, 281.6377, 281.5696, 
    281.5015, 281.4333, 281.3652, 281.2971, 281.2292, 281.1611, 281.093, 
    281.0249, 281.0085, 280.9976, 280.9871, 280.9768, 280.9666, 280.9563, 
    280.946, 280.936, 280.9258, 280.9155, 280.9053, 280.895, 280.8848, 
    280.8745, 280.8682, 280.8677, 280.8782, 280.8887, 280.8992, 280.9097, 
    280.9202, 280.9307, 280.9412, 280.9517, 280.9622, 280.9727, 280.9832, 
    280.9895, 280.968, 280.9119, 280.8557, 280.7998, 280.7437, 280.6875, 
    280.6316, 280.5754, 280.5195, 280.4634, 280.4072, 280.3513, 280.2952, 
    280.2339, 280.1646, 280.0991, 280.0337, 279.9685, 279.9031, 279.8376, 
    279.7722, 279.7068, 279.6414, 279.5759, 279.5107, 279.4453, 279.3799, 
    279.363, 279.436, 279.509, 279.5818, 279.6548, 279.7278, 279.8008, 
    279.8735, 279.9465, 280.0195, 280.0925, 280.1653, 280.2383, 280.3103, 
    280.2668, 280.1467, 280.0266, 279.9065, 279.7864, 279.6663, 279.5461, 
    279.426, 279.3059, 279.1858, 279.0654, 278.9453, 278.8252, 278.7268, 
    278.6877, 278.6855, 278.6831, 278.6809, 278.6785, 278.6763,
  276.4495, 276.4495, 276.4551, 276.4712, 276.4873, 276.5034, 276.5198, 
    276.5359, 276.552, 276.5681, 276.5845, 276.6006, 276.6243, 276.6619, 
    276.6997, 276.7375, 276.803, 276.9006, 276.9985, 277.0964, 277.1941, 
    277.292, 277.3899, 277.4878, 277.5854, 277.6833, 277.7808, 277.8782, 
    277.9756, 278.073, 278.1472, 278.2039, 278.2603, 278.3169, 278.3733, 
    278.4299, 278.4863, 278.543, 278.5994, 278.6541, 278.7078, 278.7615, 
    278.8152, 278.8689, 278.9465, 279.0354, 279.1243, 279.2131, 279.302, 
    279.3909, 279.48, 279.5688, 279.6655, 279.7776, 279.8894, 280.0015, 
    280.1133, 280.2253, 280.4031, 280.5981, 280.7932, 280.9883, 281.1833, 
    281.3784, 281.5735, 281.7686, 281.9675, 282.1667, 282.366, 282.5649, 
    282.7642, 282.9634, 283.0283, 283.0786, 283.1289, 283.1794, 283.2297, 
    283.2803, 283.3306, 283.3083, 283.2517, 283.1951, 283.1384, 283.0818, 
    283.0251, 282.9678, 282.8591, 282.7502, 282.6414, 282.5325, 282.4236, 
    282.3147, 282.2229, 282.1628, 282.103, 282.043, 281.9832, 281.9231, 
    281.8633, 281.8105, 281.8074, 281.8042, 281.8008, 281.7976, 281.7944, 
    281.791, 281.7783, 281.7654, 281.7527, 281.7397, 281.7271, 281.7141, 
    281.7014, 281.6863, 281.6636, 281.6409, 281.6182, 281.5955, 281.573, 
    281.5735, 281.5847, 281.5962, 281.6077, 281.6189, 281.6304, 281.6416, 
    281.6531, 281.6799, 281.7361, 281.792, 281.8481, 281.9041, 281.9607, 
    282.0183, 282.0759, 282.1338, 282.1914, 282.249, 282.3066, 282.3643, 
    282.4221, 282.4768, 282.5283, 282.5796, 282.6311, 282.6824, 282.7188, 
    282.7551, 282.7915, 282.8279, 282.8643, 282.9006, 282.9373, 282.9736, 
    283.01, 283.033, 283.0461, 283.0591, 283.0723, 283.0608, 283.0378, 
    283.0149, 282.9917, 282.9688, 282.9458, 282.9229, 282.8999, 282.8767, 
    282.8538, 282.7974, 282.7251, 282.6531, 282.585, 282.5247, 282.4644, 
    282.4041, 282.3438, 282.2834, 282.2231, 282.1628, 282.1025, 282.0425, 
    281.9822, 281.9185, 281.8542, 281.7898, 281.7283, 281.6665, 281.6047, 
    281.5432, 281.4814, 281.4197, 281.3579, 281.2964, 281.2346, 281.1729, 
    281.1113, 281.0916, 281.0762, 281.0618, 281.0476, 281.0334, 281.0193, 
    281.0051, 280.991, 280.9768, 280.9626, 280.9485, 280.9343, 280.9202, 
    280.906, 280.895, 280.8933, 280.9089, 280.9248, 280.9404, 280.9563, 
    280.9719, 280.9875, 281.0034, 281.019, 281.0347, 281.0505, 281.0662, 
    281.0786, 281.0679, 281.0024, 280.9373, 280.8718, 280.8066, 280.7412, 
    280.676, 280.6106, 280.5454, 280.48, 280.4148, 280.3494, 280.2842, 
    280.2146, 280.145, 280.0818, 280.0183, 279.9551, 279.8916, 279.8284, 
    279.7649, 279.7017, 279.6384, 279.575, 279.5117, 279.4482, 279.385, 
    279.3691, 279.4414, 279.5137, 279.5859, 279.6582, 279.7305, 279.8027, 
    279.875, 279.9473, 280.0195, 280.0918, 280.1641, 280.2363, 280.3071, 
    280.2461, 280.1228, 279.9995, 279.8762, 279.7529, 279.6296, 279.5063, 
    279.3831, 279.2598, 279.1365, 279.0132, 278.8901, 278.7668, 278.6775, 
    278.6445, 278.6414, 278.6379, 278.6348, 278.6313, 278.6282,
  276.4971, 276.5029, 276.5132, 276.5317, 276.55, 276.5684, 276.5869, 
    276.6052, 276.6238, 276.6421, 276.6604, 276.679, 276.7075, 276.7556, 
    276.8035, 276.8516, 276.9207, 277.0149, 277.1089, 277.2031, 277.2971, 
    277.3914, 277.4856, 277.5796, 277.6738, 277.7678, 277.8616, 277.9551, 
    278.0486, 278.1423, 278.218, 278.2803, 278.3423, 278.4045, 278.4666, 
    278.5288, 278.5911, 278.6531, 278.7153, 278.7749, 278.833, 278.8914, 
    278.9497, 279.0081, 279.0847, 279.1699, 279.2554, 279.3408, 279.426, 
    279.5115, 279.5967, 279.6821, 279.7783, 279.8953, 280.012, 280.1289, 
    280.2456, 280.3625, 280.53, 280.7107, 280.8914, 281.072, 281.2527, 
    281.4336, 281.6143, 281.7949, 281.9812, 282.1675, 282.354, 282.5403, 
    282.7266, 282.9128, 282.9958, 283.0679, 283.1399, 283.2119, 283.2839, 
    283.356, 283.428, 283.4006, 283.3262, 283.2517, 283.1772, 283.103, 
    283.0286, 282.9536, 282.8389, 282.7244, 282.6099, 282.4954, 282.3806, 
    282.2661, 282.1748, 282.1272, 282.0796, 282.032, 281.9844, 281.9368, 
    281.8892, 281.8472, 281.843, 281.8391, 281.835, 281.8311, 281.8269, 
    281.8228, 281.8057, 281.7883, 281.7712, 281.7542, 281.7368, 281.7197, 
    281.7024, 281.6836, 281.6587, 281.634, 281.6094, 281.5845, 281.5598, 
    281.5667, 281.5886, 281.6104, 281.6323, 281.6541, 281.676, 281.6978, 
    281.7197, 281.7534, 281.8096, 281.8657, 281.9219, 281.978, 282.0349, 
    282.0935, 282.1519, 282.2102, 282.2686, 282.3269, 282.3853, 282.4436, 
    282.5022, 282.5583, 282.6118, 282.6655, 282.719, 282.7725, 282.8054, 
    282.8384, 282.8716, 282.9045, 282.9375, 282.9705, 283.0037, 283.0366, 
    283.0696, 283.0923, 283.1074, 283.1226, 283.1377, 283.1191, 283.085, 
    283.0508, 283.0164, 282.9822, 282.948, 282.9136, 282.8794, 282.845, 
    282.8108, 282.7507, 282.6787, 282.6067, 282.5403, 282.4846, 282.4287, 
    282.3728, 282.3171, 282.2612, 282.2053, 282.1497, 282.0938, 282.0378, 
    281.9822, 281.9238, 281.8647, 281.8059, 281.7507, 281.6953, 281.6401, 
    281.5847, 281.5293, 281.4741, 281.4187, 281.3635, 281.3081, 281.2529, 
    281.1975, 281.1746, 281.1548, 281.1362, 281.1182, 281.1001, 281.082, 
    281.064, 281.0459, 281.0278, 281.0098, 280.9917, 280.9736, 280.9556, 
    280.9375, 280.9219, 280.9189, 280.9399, 280.9609, 280.9817, 281.0027, 
    281.0237, 281.0447, 281.0654, 281.0864, 281.1074, 281.1282, 281.1492, 
    281.1677, 281.1677, 281.093, 281.0186, 280.9441, 280.8694, 280.7949, 
    280.7205, 280.6458, 280.5713, 280.4968, 280.4221, 280.3477, 280.2732, 
    280.1953, 280.1255, 280.0642, 280.0029, 279.9417, 279.8804, 279.8191, 
    279.7578, 279.6965, 279.6353, 279.574, 279.5127, 279.4514, 279.3901, 
    279.3752, 279.447, 279.5186, 279.5901, 279.6616, 279.7332, 279.8047, 
    279.8762, 279.9478, 280.0195, 280.0911, 280.1626, 280.2341, 280.3037, 
    280.2251, 280.0989, 279.9724, 279.8459, 279.7195, 279.593, 279.4668, 
    279.3403, 279.2139, 279.0874, 278.9612, 278.8347, 278.7083, 278.6284, 
    278.6013, 278.5972, 278.5928, 278.5884, 278.5842, 278.5798,
  276.5447, 276.5566, 276.5715, 276.5923, 276.6128, 276.6335, 276.6541, 
    276.6748, 276.6953, 276.7161, 276.7366, 276.7571, 276.7908, 276.8491, 
    276.9072, 276.9656, 277.0386, 277.1289, 277.2195, 277.3098, 277.4001, 
    277.4907, 277.5811, 277.6716, 277.762, 277.8525, 277.9421, 278.032, 
    278.1216, 278.2114, 278.2888, 278.3564, 278.4243, 278.4922, 278.5601, 
    278.6277, 278.6956, 278.7634, 278.8311, 278.8955, 278.9585, 279.0215, 
    279.0842, 279.1472, 279.2229, 279.3047, 279.3865, 279.4683, 279.55, 
    279.6318, 279.7136, 279.7954, 279.8909, 280.0127, 280.1345, 280.2563, 
    280.3782, 280.4998, 280.657, 280.8232, 280.9895, 281.156, 281.3223, 
    281.4888, 281.655, 281.8215, 281.9949, 282.1685, 282.3418, 282.5154, 
    282.6887, 282.8623, 282.9636, 283.0574, 283.1509, 283.2446, 283.3381, 
    283.4319, 283.5256, 283.4929, 283.4006, 283.3086, 283.2163, 283.124, 
    283.0317, 282.9392, 282.8188, 282.6987, 282.5784, 282.458, 282.3379, 
    282.2175, 282.1267, 282.0916, 282.0562, 282.021, 281.9856, 281.9504, 
    281.915, 281.8838, 281.8789, 281.874, 281.8691, 281.8643, 281.8594, 
    281.8545, 281.8328, 281.8113, 281.7898, 281.7683, 281.7466, 281.7251, 
    281.7036, 281.6809, 281.6541, 281.6272, 281.6003, 281.5735, 281.5466, 
    281.5601, 281.5923, 281.6248, 281.657, 281.6895, 281.7217, 281.7539, 
    281.7864, 281.8269, 281.8833, 281.9395, 281.9958, 282.052, 282.1094, 
    282.1685, 282.2275, 282.2866, 282.3457, 282.4048, 282.4639, 282.5229, 
    282.5823, 282.6396, 282.6956, 282.7512, 282.8071, 282.8625, 282.8921, 
    282.9219, 282.9514, 282.981, 283.0107, 283.0403, 283.0701, 283.0996, 
    283.1294, 283.1519, 283.1689, 283.186, 283.2031, 283.1777, 283.1321, 
    283.0867, 283.041, 282.9956, 282.95, 282.9043, 282.8589, 282.8132, 
    282.7678, 282.7043, 282.6323, 282.5605, 282.4956, 282.4443, 282.3931, 
    282.3416, 282.2903, 282.239, 282.1875, 282.1362, 282.0847, 282.0334, 
    281.9822, 281.929, 281.8755, 281.822, 281.7732, 281.7241, 281.6753, 
    281.6262, 281.5774, 281.5286, 281.4795, 281.4307, 281.3818, 281.3328, 
    281.2839, 281.2576, 281.2334, 281.2109, 281.189, 281.1667, 281.1448, 
    281.1228, 281.1008, 281.0789, 281.0569, 281.0349, 281.0129, 280.991, 
    280.969, 280.9487, 280.9446, 280.9707, 280.9968, 281.0229, 281.0493, 
    281.0754, 281.1016, 281.1277, 281.1538, 281.1799, 281.2061, 281.2322, 
    281.2566, 281.2676, 281.1838, 281.0999, 281.0161, 280.9324, 280.8486, 
    280.7649, 280.6809, 280.5972, 280.5134, 280.4297, 280.3459, 280.262, 
    280.176, 280.106, 280.0466, 279.9875, 279.9282, 279.8691, 279.8098, 
    279.7505, 279.6914, 279.6321, 279.5728, 279.5137, 279.4543, 279.395, 
    279.3816, 279.4524, 279.5232, 279.5942, 279.665, 279.7358, 279.8066, 
    279.8777, 279.9485, 280.0193, 280.0903, 280.1611, 280.2319, 280.3005, 
    280.2043, 280.0747, 279.9453, 279.8157, 279.686, 279.5566, 279.427, 
    279.2974, 279.168, 279.0383, 278.9089, 278.7793, 278.6497, 278.5793, 
    278.5581, 278.553, 278.5476, 278.5422, 278.5369, 278.5317,
  276.5923, 276.6101, 276.6299, 276.6526, 276.6755, 276.6985, 276.7212, 
    276.7441, 276.7671, 276.7898, 276.8127, 276.8354, 276.874, 276.9426, 
    277.011, 277.0796, 277.1562, 277.2429, 277.3298, 277.4165, 277.5032, 
    277.5901, 277.6768, 277.7634, 277.8503, 277.937, 278.0229, 278.1089, 
    278.1948, 278.2805, 278.3594, 278.4329, 278.5063, 278.5798, 278.6533, 
    278.7266, 278.8, 278.8735, 278.947, 279.0164, 279.084, 279.1514, 279.219, 
    279.2864, 279.3611, 279.4395, 279.5176, 279.5957, 279.6741, 279.7522, 
    279.8306, 279.9087, 280.0037, 280.1304, 280.2571, 280.3838, 280.5105, 
    280.6372, 280.7839, 280.9358, 281.0879, 281.24, 281.3918, 281.5439, 
    281.696, 281.8481, 282.0085, 282.1692, 282.3298, 282.4905, 282.6511, 
    282.8115, 282.9314, 283.0466, 283.1619, 283.2771, 283.3923, 283.5078, 
    283.623, 283.5852, 283.4751, 283.3652, 283.2551, 283.145, 283.0352, 
    282.9248, 282.7988, 282.6729, 282.5469, 282.4209, 282.2949, 282.1689, 
    282.0786, 282.0557, 282.033, 282.01, 281.9871, 281.9641, 281.9412, 
    281.9204, 281.9146, 281.9089, 281.9033, 281.8977, 281.8921, 281.886, 
    281.8601, 281.8342, 281.8083, 281.7825, 281.7566, 281.7307, 281.7046, 
    281.678, 281.6492, 281.6204, 281.5913, 281.5625, 281.5334, 281.5535, 
    281.5962, 281.6389, 281.6819, 281.7246, 281.7673, 281.8101, 281.853, 
    281.9004, 281.9568, 282.0132, 282.0696, 282.126, 282.1836, 282.2434, 
    282.3032, 282.363, 282.4229, 282.4827, 282.5425, 282.6025, 282.6624, 
    282.7212, 282.7791, 282.8372, 282.895, 282.9526, 282.9788, 283.0051, 
    283.0312, 283.0576, 283.084, 283.1101, 283.1365, 283.1626, 283.189, 
    283.2112, 283.2302, 283.2495, 283.2686, 283.2361, 283.1792, 283.1226, 
    283.0657, 283.0088, 282.9519, 282.8953, 282.8384, 282.7815, 282.7249, 
    282.6577, 282.5859, 282.5142, 282.4509, 282.4041, 282.3572, 282.3103, 
    282.2634, 282.2166, 282.1697, 282.1228, 282.0759, 282.0291, 281.9822, 
    281.9343, 281.8862, 281.8381, 281.7957, 281.7529, 281.7104, 281.668, 
    281.6255, 281.583, 281.5403, 281.4978, 281.4553, 281.4128, 281.3704, 
    281.3406, 281.312, 281.2854, 281.2595, 281.2336, 281.2078, 281.1819, 
    281.156, 281.1299, 281.104, 281.0781, 281.0522, 281.0264, 281.0005, 
    280.9756, 280.9702, 281.0017, 281.033, 281.0645, 281.0957, 281.1272, 
    281.1584, 281.1899, 281.2212, 281.2527, 281.2839, 281.3154, 281.3457, 
    281.3674, 281.2744, 281.1814, 281.0884, 280.9954, 280.9023, 280.8091, 
    280.7161, 280.623, 280.53, 280.437, 280.344, 280.251, 280.1567, 280.0864, 
    280.0293, 279.9722, 279.9148, 279.8577, 279.8005, 279.7434, 279.686, 
    279.6289, 279.5718, 279.5146, 279.4573, 279.4001, 279.3877, 279.4578, 
    279.5281, 279.5981, 279.6685, 279.7385, 279.8088, 279.8789, 279.9492, 
    280.0193, 280.0896, 280.1597, 280.23, 280.2974, 280.1836, 280.0508, 
    279.9182, 279.7854, 279.6528, 279.52, 279.3875, 279.2546, 279.1221, 
    278.9893, 278.8567, 278.7239, 278.5913, 278.5303, 278.5149, 278.5088, 
    278.5024, 278.4961, 278.4897, 278.4834,
  276.6399, 276.6638, 276.6882, 276.7131, 276.7383, 276.7634, 276.7886, 
    276.8135, 276.8386, 276.8638, 276.8887, 276.9138, 276.9573, 277.0361, 
    277.1147, 277.1934, 277.2742, 277.3572, 277.4402, 277.5232, 277.6062, 
    277.6892, 277.7725, 277.8555, 277.9385, 278.0215, 278.1035, 278.1855, 
    278.2678, 278.3499, 278.4302, 278.5093, 278.5884, 278.6675, 278.7466, 
    278.8257, 278.9048, 278.9839, 279.0627, 279.1372, 279.2092, 279.2815, 
    279.3535, 279.4255, 279.4995, 279.574, 279.6487, 279.7234, 279.7981, 
    279.8728, 279.9473, 280.022, 280.1162, 280.2478, 280.3796, 280.5112, 
    280.6428, 280.7744, 280.9106, 281.0483, 281.186, 281.3237, 281.4614, 
    281.5991, 281.7368, 281.8745, 282.0222, 282.1702, 282.3179, 282.4656, 
    282.6133, 282.761, 282.8989, 283.0359, 283.1729, 283.3098, 283.4465, 
    283.5835, 283.7205, 283.6775, 283.5498, 283.4219, 283.2939, 283.1663, 
    283.0383, 282.9104, 282.7788, 282.6472, 282.5154, 282.3838, 282.2522, 
    282.1204, 282.0308, 282.02, 282.0095, 281.9988, 281.9883, 281.9775, 
    281.967, 281.9568, 281.9504, 281.9438, 281.9375, 281.9309, 281.9246, 
    281.9177, 281.8875, 281.8572, 281.8269, 281.7966, 281.7664, 281.7361, 
    281.7058, 281.6753, 281.6443, 281.6135, 281.5825, 281.5515, 281.5205, 
    281.5466, 281.6001, 281.6533, 281.7065, 281.7598, 281.813, 281.8662, 
    281.9194, 281.9739, 282.0305, 282.0869, 282.1433, 282.2, 282.2578, 
    282.3184, 282.3789, 282.4395, 282.5, 282.5605, 282.6213, 282.6819, 
    282.7424, 282.8027, 282.8628, 282.9229, 282.9832, 283.0427, 283.0654, 
    283.0884, 283.1113, 283.1343, 283.157, 283.1799, 283.2029, 283.2258, 
    283.2485, 283.2705, 283.2917, 283.313, 283.3342, 283.2944, 283.2263, 
    283.1584, 283.0903, 283.0222, 282.9541, 282.886, 282.8179, 282.7498, 
    282.6816, 282.6111, 282.5396, 282.4678, 282.4062, 282.364, 282.3215, 
    282.2791, 282.2366, 282.1943, 282.1519, 282.1094, 282.0669, 282.0247, 
    281.9822, 281.9395, 281.8967, 281.8542, 281.8181, 281.782, 281.7456, 
    281.7095, 281.6733, 281.6372, 281.6011, 281.5649, 281.5288, 281.4927, 
    281.4565, 281.4236, 281.3909, 281.3601, 281.3301, 281.3003, 281.2705, 
    281.2407, 281.2109, 281.1812, 281.1511, 281.1213, 281.0916, 281.0618, 
    281.032, 281.0024, 280.9958, 281.0325, 281.0691, 281.1057, 281.1423, 
    281.1787, 281.2153, 281.252, 281.2886, 281.3252, 281.3618, 281.3984, 
    281.4348, 281.4673, 281.365, 281.2627, 281.1604, 281.0581, 280.9558, 
    280.8535, 280.7512, 280.6492, 280.5469, 280.4446, 280.3423, 280.24, 
    280.1375, 280.0669, 280.0117, 279.9565, 279.9016, 279.8464, 279.7913, 
    279.7361, 279.6809, 279.6257, 279.5706, 279.5156, 279.4604, 279.4053, 
    279.3938, 279.4634, 279.5327, 279.6023, 279.6719, 279.7412, 279.8108, 
    279.8804, 279.9497, 280.0193, 280.0889, 280.1582, 280.2278, 280.2939, 
    280.1626, 280.0269, 279.8911, 279.7551, 279.6194, 279.4834, 279.3477, 
    279.2119, 279.0759, 278.9402, 278.8044, 278.6685, 278.5327, 278.4812, 
    278.4717, 278.4646, 278.4573, 278.45, 278.4426, 278.4353,
  276.6992, 276.728, 276.7566, 276.7852, 276.814, 276.8425, 276.8711, 
    276.8999, 276.9285, 276.957, 276.9856, 277.0144, 277.0637, 277.1531, 
    277.2424, 277.3315, 277.4209, 277.5103, 277.5994, 277.6887, 277.7778, 
    277.8672, 277.9565, 278.0457, 278.135, 278.2241, 278.2961, 278.3682, 
    278.4404, 278.5125, 278.5847, 278.6567, 278.7288, 278.801, 278.873, 
    278.9453, 279.0173, 279.0894, 279.1616, 279.2341, 279.3069, 279.3796, 
    279.4524, 279.5251, 279.5979, 279.6709, 279.7437, 279.8164, 279.8892, 
    279.9619, 280.0347, 280.1074, 280.2009, 280.3337, 280.4663, 280.5991, 
    280.7319, 280.8645, 280.9973, 281.1301, 281.2627, 281.3955, 281.5283, 
    281.6609, 281.7937, 281.9263, 282.0574, 282.1882, 282.3193, 282.4502, 
    282.5813, 282.7122, 282.843, 282.9741, 283.105, 283.2361, 283.3669, 
    283.4978, 283.6289, 283.5889, 283.4678, 283.3469, 283.2258, 283.105, 
    282.9839, 282.863, 282.7419, 282.6211, 282.5, 282.3792, 282.2583, 
    282.1372, 282.0562, 282.0503, 282.0444, 282.0386, 282.0327, 282.0269, 
    282.021, 282.0149, 282.009, 282.0032, 281.9973, 281.9915, 281.9856, 
    281.9795, 281.9504, 281.9214, 281.8923, 281.8633, 281.8342, 281.8052, 
    281.7761, 281.7471, 281.718, 281.6892, 281.6602, 281.6311, 281.6021, 
    281.6201, 281.6606, 281.7014, 281.7419, 281.7825, 281.823, 281.8635, 
    281.9041, 281.9446, 281.9851, 282.0256, 282.0662, 282.1067, 282.1562, 
    282.2229, 282.2893, 282.356, 282.4226, 282.4893, 282.5559, 282.6226, 
    282.6892, 282.7559, 282.8223, 282.8889, 282.9556, 283.0217, 283.051, 
    283.0801, 283.1094, 283.1384, 283.1677, 283.197, 283.2261, 283.2554, 
    283.2844, 283.3137, 283.343, 283.3721, 283.4014, 283.3589, 283.283, 
    283.2073, 283.1313, 283.0554, 282.9795, 282.9036, 282.8276, 282.7517, 
    282.676, 282.6001, 282.5242, 282.4482, 282.3855, 282.3472, 282.3088, 
    282.2708, 282.2324, 282.1941, 282.156, 282.1177, 282.0793, 282.041, 
    282.0029, 281.9646, 281.9263, 281.8882, 281.855, 281.8215, 281.7883, 
    281.7551, 281.7217, 281.6885, 281.655, 281.6218, 281.5886, 281.5552, 
    281.522, 281.4888, 281.4553, 281.4209, 281.386, 281.3511, 281.3162, 
    281.2812, 281.2461, 281.2112, 281.1763, 281.1414, 281.1064, 281.0715, 
    281.0364, 281.0015, 280.9895, 281.02, 281.0505, 281.0813, 281.1118, 
    281.1426, 281.1731, 281.2036, 281.2344, 281.2649, 281.2954, 281.3262, 
    281.3567, 281.3853, 281.2898, 281.1943, 281.0989, 281.0034, 280.9077, 
    280.8123, 280.7168, 280.6213, 280.5259, 280.4304, 280.335, 280.2393, 
    280.1438, 280.0774, 280.0242, 279.9709, 279.9177, 279.8645, 279.8113, 
    279.7581, 279.7048, 279.6516, 279.5984, 279.5452, 279.4919, 279.4387, 
    279.425, 279.4844, 279.5439, 279.6033, 279.6626, 279.7222, 279.7815, 
    279.8411, 279.9004, 279.96, 280.0193, 280.0786, 280.1382, 280.1946, 
    280.0728, 279.9509, 279.8293, 279.7075, 279.5857, 279.4641, 279.3423, 
    279.2205, 279.0989, 278.9771, 278.8552, 278.7336, 278.6118, 278.5671, 
    278.5581, 278.5491, 278.5403, 278.5312, 278.5222, 278.5132,
  276.7642, 276.7969, 276.8298, 276.8625, 276.8953, 276.9282, 276.9609, 
    276.9937, 277.0266, 277.0593, 277.0923, 277.125, 277.1809, 277.281, 
    277.3809, 277.481, 277.5811, 277.6809, 277.781, 277.8811, 277.981, 
    278.0811, 278.1812, 278.281, 278.3811, 278.4807, 278.54, 278.5994, 
    278.6587, 278.718, 278.7773, 278.8369, 278.8962, 278.9556, 279.0149, 
    279.0742, 279.1335, 279.1929, 279.2524, 279.3201, 279.3918, 279.4634, 
    279.5352, 279.6067, 279.6785, 279.75, 279.8218, 279.8936, 279.9651, 
    280.0369, 280.1084, 280.1802, 280.2727, 280.4048, 280.5369, 280.6689, 
    280.801, 280.9331, 281.0654, 281.1975, 281.3296, 281.4617, 281.5938, 
    281.7258, 281.8579, 281.9897, 282.1021, 282.2146, 282.3269, 282.4392, 
    282.5518, 282.6641, 282.7764, 282.8887, 283.0012, 283.1135, 283.2258, 
    283.3381, 283.4507, 283.417, 283.3142, 283.2114, 283.1086, 283.0059, 
    282.9031, 282.8005, 282.6978, 282.595, 282.4922, 282.3894, 282.2866, 
    282.1838, 282.1152, 282.1106, 282.106, 282.1013, 282.0967, 282.0923, 
    282.0876, 282.083, 282.0784, 282.0737, 282.0691, 282.0647, 282.0601, 
    282.0552, 282.0298, 282.0046, 281.9795, 281.9541, 281.929, 281.9036, 
    281.8784, 281.8533, 281.8279, 281.8027, 281.7773, 281.7522, 281.7268, 
    281.7305, 281.7476, 281.7649, 281.782, 281.7991, 281.8164, 281.8335, 
    281.8506, 281.8679, 281.885, 281.9021, 281.9194, 281.9365, 281.9739, 
    282.0488, 282.124, 282.1992, 282.2742, 282.3494, 282.4246, 282.4998, 
    282.5747, 282.6499, 282.7251, 282.8, 282.8752, 282.95, 282.9897, 
    283.0298, 283.0698, 283.1096, 283.1497, 283.1897, 283.2295, 283.2695, 
    283.3096, 283.3494, 283.3894, 283.4294, 283.4692, 283.426, 283.344, 
    283.262, 283.1799, 283.0977, 283.0156, 282.9336, 282.8513, 282.7693, 
    282.6873, 282.6052, 282.5229, 282.4409, 282.3755, 282.3413, 282.3069, 
    282.2727, 282.2385, 282.2043, 282.1702, 282.1357, 282.1016, 282.0674, 
    282.0332, 281.9988, 281.9646, 281.9304, 281.8984, 281.8662, 281.8342, 
    281.8022, 281.77, 281.738, 281.7061, 281.6741, 281.6418, 281.6099, 
    281.5779, 281.5457, 281.5137, 281.4758, 281.4351, 281.3945, 281.3538, 
    281.3132, 281.2725, 281.2319, 281.1912, 281.1506, 281.1099, 281.0693, 
    281.0286, 280.988, 280.9683, 280.9878, 281.0073, 281.0269, 281.0461, 
    281.0657, 281.0852, 281.1047, 281.124, 281.1436, 281.1631, 281.1826, 
    281.2019, 281.22, 281.1384, 281.0571, 280.9758, 280.8945, 280.813, 
    280.7317, 280.6504, 280.5691, 280.4875, 280.4062, 280.325, 280.2437, 
    280.1621, 280.1013, 280.05, 279.9988, 279.9473, 279.896, 279.8447, 
    279.7935, 279.7419, 279.6907, 279.6394, 279.5881, 279.5366, 279.4854, 
    279.4678, 279.5127, 279.5579, 279.603, 279.6479, 279.6931, 279.738, 
    279.7832, 279.8281, 279.8733, 279.9182, 279.9634, 280.0083, 280.051, 
    279.9512, 279.8513, 279.7517, 279.6519, 279.5522, 279.4524, 279.3525, 
    279.2529, 279.1531, 279.0535, 278.9536, 278.8538, 278.7542, 278.7151, 
    278.7041, 278.6929, 278.6819, 278.6709, 278.6599, 278.6489,
  276.8289, 276.866, 276.9028, 276.9399, 276.9768, 277.0137, 277.0508, 
    277.0876, 277.1248, 277.1616, 277.1987, 277.2356, 277.2981, 277.4087, 
    277.5195, 277.6304, 277.741, 277.8518, 277.9626, 278.0735, 278.1841, 
    278.2949, 278.4058, 278.5164, 278.6272, 278.7373, 278.7839, 278.8306, 
    278.8772, 278.9236, 278.9702, 279.0168, 279.0635, 279.1101, 279.1567, 
    279.2034, 279.25, 279.2966, 279.3433, 279.406, 279.4766, 279.5471, 
    279.6177, 279.6882, 279.7588, 279.8293, 279.8999, 279.9707, 280.0413, 
    280.1118, 280.1824, 280.2529, 280.3445, 280.4758, 280.6074, 280.7388, 
    280.8704, 281.002, 281.1333, 281.2649, 281.3962, 281.5278, 281.6592, 
    281.7908, 281.9221, 282.0532, 282.147, 282.2407, 282.3345, 282.4282, 
    282.5222, 282.616, 282.7097, 282.8035, 282.8972, 282.991, 283.0847, 
    283.1785, 283.2722, 283.2451, 283.1604, 283.0759, 282.9915, 282.907, 
    282.8223, 282.7378, 282.6533, 282.5688, 282.4844, 282.3997, 282.3152, 
    282.2307, 282.1743, 282.1709, 282.1675, 282.1643, 282.1609, 282.1577, 
    282.1543, 282.1509, 282.1477, 282.1443, 282.1409, 282.1377, 282.1343, 
    282.1309, 282.1094, 282.0879, 282.0664, 282.0449, 282.0234, 282.002, 
    281.9807, 281.9592, 281.9377, 281.9163, 281.8948, 281.8733, 281.8518, 
    281.8408, 281.8345, 281.8284, 281.8223, 281.8159, 281.8098, 281.8035, 
    281.7974, 281.7913, 281.7849, 281.7788, 281.7727, 281.7664, 281.7913, 
    281.875, 281.9587, 282.0422, 282.126, 282.2095, 282.2932, 282.3767, 
    282.4604, 282.5439, 282.6277, 282.7112, 282.7949, 282.8782, 282.9287, 
    282.9795, 283.0303, 283.0808, 283.1316, 283.1824, 283.2329, 283.2837, 
    283.3345, 283.3853, 283.4358, 283.4866, 283.5374, 283.4934, 283.405, 
    283.3167, 283.2283, 283.1401, 283.0518, 282.9634, 282.8752, 282.7869, 
    282.6985, 282.6101, 282.522, 282.4336, 282.3655, 282.3352, 282.3049, 
    282.2749, 282.2446, 282.2144, 282.1841, 282.1541, 282.1238, 282.0935, 
    282.0632, 282.0332, 282.0029, 281.9727, 281.9419, 281.9111, 281.8801, 
    281.8494, 281.8186, 281.7876, 281.7568, 281.7261, 281.6953, 281.6643, 
    281.6335, 281.6028, 281.5718, 281.5305, 281.4841, 281.4377, 281.3916, 
    281.3452, 281.2988, 281.2524, 281.2061, 281.1599, 281.1135, 281.0671, 
    281.0208, 280.9744, 280.9473, 280.9556, 280.9639, 280.9722, 280.9807, 
    280.989, 280.9973, 281.0056, 281.0139, 281.0222, 281.0308, 281.0391, 
    281.0474, 281.0544, 280.9873, 280.9199, 280.8528, 280.7856, 280.7183, 
    280.6511, 280.584, 280.5166, 280.4495, 280.3821, 280.3149, 280.2478, 
    280.1804, 280.1255, 280.0759, 280.0266, 279.9771, 279.9275, 279.8782, 
    279.8286, 279.7793, 279.7297, 279.6804, 279.6309, 279.5813, 279.532, 
    279.5105, 279.5413, 279.5718, 279.6025, 279.6333, 279.6638, 279.6946, 
    279.7251, 279.7559, 279.7866, 279.8171, 279.8479, 279.8787, 279.9075, 
    279.8296, 279.7517, 279.6741, 279.5962, 279.5186, 279.4407, 279.363, 
    279.2852, 279.2075, 279.1296, 279.052, 278.9741, 278.8962, 278.8628, 
    278.8499, 278.8367, 278.8237, 278.8108, 278.7976, 278.7847,
  276.8938, 276.9348, 276.9761, 277.0171, 277.0583, 277.0994, 277.1406, 
    277.1816, 277.2229, 277.2639, 277.3052, 277.3462, 277.415, 277.5366, 
    277.6582, 277.7795, 277.9011, 278.0227, 278.1443, 278.2656, 278.3872, 
    278.5088, 278.6304, 278.7517, 278.8733, 278.9939, 279.0278, 279.0615, 
    279.0955, 279.1294, 279.1631, 279.197, 279.231, 279.2646, 279.2986, 
    279.3325, 279.3662, 279.4001, 279.4341, 279.4919, 279.5615, 279.6309, 
    279.7004, 279.7698, 279.8394, 279.9087, 279.9783, 280.0476, 280.1172, 
    280.1865, 280.2561, 280.3254, 280.4163, 280.5471, 280.678, 280.8088, 
    280.9397, 281.0706, 281.2014, 281.3323, 281.4631, 281.594, 281.7249, 
    281.8555, 281.9863, 282.1167, 282.1919, 282.2671, 282.3423, 282.4175, 
    282.4927, 282.5679, 282.6428, 282.718, 282.7932, 282.8684, 282.9436, 
    283.0188, 283.094, 283.0732, 283.0068, 282.9404, 282.8743, 282.8079, 
    282.7417, 282.6753, 282.6089, 282.5427, 282.4763, 282.4099, 282.3438, 
    282.2773, 282.2334, 282.2312, 282.2292, 282.2271, 282.2251, 282.2231, 
    282.2209, 282.219, 282.2168, 282.2148, 282.2129, 282.2107, 282.2087, 
    282.2063, 282.1887, 282.1711, 282.1533, 282.1357, 282.1182, 282.1003, 
    282.0828, 282.0652, 282.0474, 282.0298, 282.0122, 281.9944, 281.9768, 
    281.9512, 281.9214, 281.8918, 281.8623, 281.8328, 281.8032, 281.7737, 
    281.7441, 281.7146, 281.6851, 281.6555, 281.626, 281.5962, 281.6089, 
    281.7012, 281.7932, 281.8853, 281.9775, 282.0696, 282.1619, 282.2539, 
    282.3459, 282.4382, 282.5303, 282.6223, 282.7146, 282.8062, 282.8677, 
    282.9292, 282.9907, 283.052, 283.1135, 283.175, 283.2366, 283.2979, 
    283.3594, 283.4209, 283.4824, 283.5437, 283.6052, 283.5605, 283.4661, 
    283.3713, 283.2769, 283.1824, 283.0879, 282.9934, 282.8989, 282.8042, 
    282.7097, 282.6152, 282.5208, 282.4263, 282.3555, 282.3293, 282.303, 
    282.2769, 282.2507, 282.2246, 282.1982, 282.1721, 282.146, 282.1199, 
    282.0935, 282.0674, 282.0413, 282.0149, 281.9854, 281.9558, 281.926, 
    281.8965, 281.8669, 281.8374, 281.8079, 281.7781, 281.7485, 281.719, 
    281.6895, 281.6597, 281.6301, 281.5852, 281.5332, 281.4812, 281.4292, 
    281.3772, 281.3252, 281.2732, 281.2209, 281.1689, 281.1169, 281.0649, 
    281.0129, 280.9609, 280.926, 280.9233, 280.9204, 280.9177, 280.915, 
    280.9121, 280.9094, 280.9065, 280.9038, 280.9011, 280.8982, 280.8955, 
    280.8926, 280.8892, 280.8359, 280.783, 280.7297, 280.6768, 280.6235, 
    280.5706, 280.5173, 280.4644, 280.4111, 280.3582, 280.3049, 280.252, 
    280.1987, 280.1494, 280.1018, 280.0542, 280.0068, 279.9592, 279.9116, 
    279.864, 279.8164, 279.7688, 279.7212, 279.6736, 279.626, 279.5786, 
    279.5532, 279.5696, 279.5859, 279.6021, 279.6184, 279.6348, 279.6511, 
    279.6672, 279.6836, 279.7, 279.7161, 279.7324, 279.7488, 279.7639, 
    279.708, 279.6523, 279.5964, 279.5408, 279.4849, 279.4292, 279.3733, 
    279.3176, 279.2617, 279.2061, 279.1501, 279.0945, 279.0386, 279.0107, 
    278.9956, 278.9805, 278.9656, 278.9504, 278.9353, 278.9204,
  276.9585, 277.0039, 277.0491, 277.0945, 277.1396, 277.1851, 277.2305, 
    277.2756, 277.321, 277.3662, 277.4116, 277.457, 277.5322, 277.6643, 
    277.7966, 277.929, 278.0613, 278.1936, 278.3259, 278.458, 278.5903, 
    278.7227, 278.855, 278.9873, 279.1194, 279.2505, 279.2717, 279.2927, 
    279.3137, 279.335, 279.356, 279.3772, 279.3982, 279.4192, 279.4404, 
    279.4614, 279.4827, 279.5037, 279.5247, 279.5779, 279.6462, 279.7146, 
    279.783, 279.8513, 279.9197, 279.988, 280.0564, 280.1248, 280.1931, 
    280.2615, 280.3298, 280.3982, 280.488, 280.6182, 280.7485, 280.8787, 
    281.0088, 281.1392, 281.2693, 281.3997, 281.5298, 281.6599, 281.7903, 
    281.9204, 282.0508, 282.1799, 282.2366, 282.2932, 282.3499, 282.4065, 
    282.4631, 282.5195, 282.5762, 282.6328, 282.6895, 282.7461, 282.8025, 
    282.8591, 282.9158, 282.9014, 282.8533, 282.8052, 282.7571, 282.709, 
    282.6609, 282.6128, 282.5647, 282.5166, 282.4685, 282.4204, 282.3723, 
    282.3242, 282.2925, 282.2915, 282.2908, 282.29, 282.2893, 282.2886, 
    282.2876, 282.2869, 282.2861, 282.2854, 282.2847, 282.2837, 282.283, 
    282.282, 282.2681, 282.2544, 282.2405, 282.2266, 282.2126, 282.1987, 
    282.1851, 282.1711, 282.1572, 282.1433, 282.1294, 282.1157, 282.1018, 
    282.0613, 282.0083, 281.9556, 281.9026, 281.8496, 281.7966, 281.7437, 
    281.6909, 281.6379, 281.585, 281.532, 281.4792, 281.4263, 281.4265, 
    281.5271, 281.6279, 281.7285, 281.8291, 281.9297, 282.0303, 282.1311, 
    282.2317, 282.3323, 282.4329, 282.5334, 282.6343, 282.7344, 282.8066, 
    282.8789, 282.9512, 283.0232, 283.0955, 283.1677, 283.24, 283.3123, 
    283.3843, 283.4565, 283.5288, 283.6011, 283.6733, 283.6277, 283.5269, 
    283.4263, 283.3254, 283.2249, 283.124, 283.0232, 282.9226, 282.8218, 
    282.7212, 282.6204, 282.5195, 282.4189, 282.3455, 282.3232, 282.3013, 
    282.2791, 282.2568, 282.2346, 282.2124, 282.1902, 282.1682, 282.146, 
    282.1238, 282.1016, 282.0793, 282.0571, 282.0288, 282.0005, 281.9722, 
    281.9436, 281.9153, 281.887, 281.8586, 281.8303, 281.8018, 281.7734, 
    281.7451, 281.7168, 281.6885, 281.6399, 281.5823, 281.5247, 281.4668, 
    281.4092, 281.3513, 281.2937, 281.2361, 281.1782, 281.1206, 281.0627, 
    281.0051, 280.9475, 280.905, 280.8911, 280.8772, 280.8633, 280.8494, 
    280.8354, 280.8215, 280.8076, 280.7937, 280.7798, 280.7659, 280.752, 
    280.738, 280.7236, 280.6848, 280.6458, 280.6067, 280.5679, 280.5288, 
    280.49, 280.4509, 280.4119, 280.373, 280.334, 280.2952, 280.2561, 
    280.217, 280.1736, 280.1279, 280.082, 280.0364, 279.9907, 279.9451, 
    279.8994, 279.8535, 279.8079, 279.7622, 279.7166, 279.6709, 279.625, 
    279.5959, 279.5979, 279.5999, 279.6018, 279.6038, 279.6055, 279.6074, 
    279.6094, 279.6113, 279.6133, 279.6152, 279.6169, 279.6189, 279.6201, 
    279.5864, 279.5527, 279.5188, 279.4851, 279.4512, 279.4175, 279.3838, 
    279.3499, 279.3162, 279.2822, 279.2485, 279.2146, 279.1809, 279.1584, 
    279.1414, 279.1243, 279.1072, 279.0901, 279.073, 279.0559,
  277.0232, 277.0728, 277.1223, 277.1716, 277.2212, 277.2708, 277.3201, 
    277.3696, 277.4192, 277.4685, 277.5181, 277.5676, 277.6492, 277.7922, 
    277.9353, 278.0784, 278.2214, 278.3645, 278.5073, 278.6504, 278.7935, 
    278.9365, 279.0796, 279.2227, 279.3657, 279.5071, 279.5154, 279.5239, 
    279.5322, 279.5405, 279.5488, 279.5571, 279.5654, 279.574, 279.5823, 
    279.5906, 279.5989, 279.6072, 279.6155, 279.6638, 279.7312, 279.7983, 
    279.8657, 279.9329, 280.0002, 280.0674, 280.1348, 280.2019, 280.2693, 
    280.3364, 280.4038, 280.4709, 280.5598, 280.6892, 280.8188, 280.9485, 
    281.0781, 281.2078, 281.3374, 281.467, 281.5964, 281.7261, 281.8557, 
    281.9854, 282.115, 282.2434, 282.2815, 282.3196, 282.3574, 282.3955, 
    282.4336, 282.4714, 282.5095, 282.5476, 282.5854, 282.6235, 282.6616, 
    282.6995, 282.7375, 282.7295, 282.6995, 282.6697, 282.6399, 282.6099, 
    282.5801, 282.55, 282.5203, 282.4905, 282.4604, 282.4307, 282.4006, 
    282.3708, 282.3516, 282.3521, 282.3525, 282.353, 282.3535, 282.354, 
    282.3545, 282.355, 282.3555, 282.356, 282.3564, 282.3569, 282.3574, 
    282.3577, 282.3477, 282.3376, 282.3274, 282.3174, 282.3074, 282.2971, 
    282.2871, 282.2771, 282.2671, 282.2568, 282.2468, 282.2368, 282.2268, 
    282.1716, 282.0952, 282.019, 281.9426, 281.8665, 281.79, 281.7139, 
    281.6375, 281.5613, 281.4849, 281.4087, 281.3325, 281.2561, 281.2441, 
    281.3533, 281.4624, 281.5715, 281.6807, 281.7898, 281.8989, 282.0081, 
    282.1172, 282.2263, 282.3354, 282.4446, 282.554, 282.6626, 282.7456, 
    282.8286, 282.9116, 282.9944, 283.0774, 283.1604, 283.2434, 283.3264, 
    283.4094, 283.4924, 283.5752, 283.6582, 283.7412, 283.6948, 283.5879, 
    283.481, 283.374, 283.2671, 283.1602, 283.0532, 282.9463, 282.8394, 
    282.7324, 282.6255, 282.5186, 282.4116, 282.3354, 282.3174, 282.2993, 
    282.281, 282.2629, 282.2449, 282.2266, 282.2085, 282.1904, 282.1721, 
    282.1541, 282.136, 282.1177, 282.0994, 282.0723, 282.0452, 282.0181, 
    281.991, 281.9639, 281.9365, 281.9094, 281.8823, 281.8552, 281.8281, 
    281.801, 281.7737, 281.7466, 281.6948, 281.6313, 281.5679, 281.5046, 
    281.4412, 281.3777, 281.3142, 281.251, 281.1875, 281.124, 281.0608, 
    280.9973, 280.9338, 280.8838, 280.8589, 280.8337, 280.8088, 280.7837, 
    280.7585, 280.7336, 280.7085, 280.6836, 280.6584, 280.6335, 280.6084, 
    280.5833, 280.5583, 280.5334, 280.5085, 280.4839, 280.459, 280.4341, 
    280.4092, 280.3845, 280.3596, 280.3347, 280.3098, 280.2852, 280.2603, 
    280.2354, 280.1975, 280.1538, 280.1099, 280.0662, 280.0222, 279.9785, 
    279.9346, 279.8909, 279.8469, 279.8032, 279.7593, 279.7156, 279.6716, 
    279.6389, 279.6262, 279.6138, 279.6013, 279.5889, 279.5764, 279.564, 
    279.5515, 279.5391, 279.5266, 279.5142, 279.5017, 279.489, 279.4766, 
    279.4648, 279.4531, 279.4412, 279.4294, 279.4177, 279.4058, 279.394, 
    279.3823, 279.3704, 279.3586, 279.3467, 279.335, 279.3232, 279.3064, 
    279.2874, 279.2681, 279.249, 279.23, 279.2109, 279.1917,
  277.0881, 277.1416, 277.1953, 277.249, 277.3027, 277.3562, 277.4099, 
    277.4636, 277.5173, 277.5708, 277.6245, 277.6782, 277.7664, 277.9202, 
    278.074, 278.2275, 278.3813, 278.5352, 278.689, 278.8428, 278.9966, 
    279.1504, 279.3042, 279.458, 279.6118, 279.7637, 279.7593, 279.7549, 
    279.7505, 279.7461, 279.7417, 279.7373, 279.7329, 279.7285, 279.7241, 
    279.7197, 279.7153, 279.7107, 279.7063, 279.7498, 279.8159, 279.8821, 
    279.9482, 280.0144, 280.0806, 280.1467, 280.2129, 280.2791, 280.3452, 
    280.4114, 280.4775, 280.5437, 280.6316, 280.7605, 280.8894, 281.0183, 
    281.1475, 281.2764, 281.4053, 281.5344, 281.6633, 281.7922, 281.9211, 
    282.0503, 282.1792, 282.3069, 282.3262, 282.3457, 282.365, 282.3845, 
    282.4041, 282.4233, 282.4429, 282.4622, 282.4817, 282.501, 282.5205, 
    282.5398, 282.5593, 282.5576, 282.5459, 282.5342, 282.5225, 282.511, 
    282.4993, 282.4875, 282.4758, 282.4641, 282.4526, 282.4409, 282.4292, 
    282.4175, 282.4104, 282.4124, 282.4141, 282.4158, 282.4175, 282.4194, 
    282.4211, 282.4229, 282.4246, 282.4263, 282.4282, 282.4299, 282.4316, 
    282.4333, 282.427, 282.4207, 282.4146, 282.4082, 282.4019, 282.3955, 
    282.3894, 282.3831, 282.3767, 282.3706, 282.3643, 282.3579, 282.3516, 
    282.282, 282.1821, 282.0825, 281.9829, 281.8833, 281.7837, 281.6838, 
    281.5842, 281.4846, 281.385, 281.2854, 281.1858, 281.0859, 281.0618, 
    281.1794, 281.2971, 281.4148, 281.5322, 281.6499, 281.7676, 281.8853, 
    282.0029, 282.1206, 282.2383, 282.356, 282.4734, 282.5908, 282.6846, 
    282.7783, 282.8721, 282.9656, 283.0593, 283.1531, 283.2468, 283.3406, 
    283.4343, 283.5281, 283.6218, 283.7156, 283.8093, 283.762, 283.6489, 
    283.5356, 283.4226, 283.3093, 283.1963, 283.083, 282.97, 282.8569, 
    282.7437, 282.6306, 282.5173, 282.4043, 282.3254, 282.3113, 282.2974, 
    282.2832, 282.269, 282.2549, 282.2407, 282.2266, 282.2124, 282.1985, 
    282.1843, 282.1702, 282.156, 282.1416, 282.1157, 282.0898, 282.064, 
    282.0381, 282.0122, 281.9863, 281.9604, 281.9343, 281.9084, 281.8826, 
    281.8567, 281.8308, 281.8049, 281.7495, 281.6804, 281.6113, 281.5422, 
    281.4731, 281.4041, 281.335, 281.2659, 281.1968, 281.1277, 281.0586, 
    280.9895, 280.9204, 280.8628, 280.8267, 280.7905, 280.7542, 280.718, 
    280.6819, 280.6458, 280.6096, 280.5735, 280.5371, 280.501, 280.4648, 
    280.4287, 280.3928, 280.3823, 280.3716, 280.3608, 280.3501, 280.3394, 
    280.3286, 280.3179, 280.3074, 280.2966, 280.2859, 280.2751, 280.2644, 
    280.2537, 280.2217, 280.1797, 280.1377, 280.0957, 280.054, 280.012, 
    279.97, 279.928, 279.886, 279.844, 279.8022, 279.7603, 279.7183, 
    279.6816, 279.6548, 279.6279, 279.6011, 279.5742, 279.5474, 279.5205, 
    279.4937, 279.4668, 279.4399, 279.4131, 279.3862, 279.3594, 279.333, 
    279.3433, 279.3535, 279.3635, 279.3738, 279.384, 279.3943, 279.4043, 
    279.4146, 279.4248, 279.4348, 279.4451, 279.4553, 279.4656, 279.4543, 
    279.4331, 279.4119, 279.3909, 279.3696, 279.3486, 279.3274,
  277.123, 277.1741, 277.2249, 277.2759, 277.3267, 277.3774, 277.4285, 
    277.4792, 277.53, 277.5811, 277.6318, 277.6829, 277.769, 277.9226, 
    278.0762, 278.2297, 278.3833, 278.5369, 278.6907, 278.8442, 278.9978, 
    279.1514, 279.3049, 279.4585, 279.6121, 279.7642, 279.7661, 279.7678, 
    279.7698, 279.7717, 279.7737, 279.7756, 279.7776, 279.7795, 279.7812, 
    279.7832, 279.7852, 279.7871, 279.7891, 279.8252, 279.8777, 279.9299, 
    279.9824, 280.0349, 280.0874, 280.1396, 280.1921, 280.2446, 280.2971, 
    280.3494, 280.4019, 280.4543, 280.5337, 280.6648, 280.7957, 280.9265, 
    281.0576, 281.1885, 281.3193, 281.4504, 281.5813, 281.7122, 281.8433, 
    281.9741, 282.105, 282.2349, 282.261, 282.2874, 282.3135, 282.3398, 
    282.366, 282.3923, 282.4187, 282.4448, 282.4712, 282.4973, 282.5237, 
    282.55, 282.5762, 282.5708, 282.55, 282.5295, 282.509, 282.4885, 282.468, 
    282.4475, 282.427, 282.4065, 282.386, 282.3655, 282.345, 282.3245, 
    282.3181, 282.3389, 282.3596, 282.3804, 282.4009, 282.4216, 282.4424, 
    282.4631, 282.4839, 282.5046, 282.5251, 282.5459, 282.5667, 282.5869, 
    282.5769, 282.5667, 282.5564, 282.5459, 282.5352, 282.5247, 282.5137, 
    282.5027, 282.4917, 282.4805, 282.469, 282.4575, 282.446, 282.3711, 
    282.2676, 282.165, 282.064, 281.9641, 281.8652, 281.7676, 281.6711, 
    281.5759, 281.4814, 281.3884, 281.2961, 281.2051, 281.1833, 281.2903, 
    281.3975, 281.5044, 281.6116, 281.7185, 281.8254, 281.9326, 282.0396, 
    282.1467, 282.2537, 282.3608, 282.4678, 282.5747, 282.6709, 282.7671, 
    282.8633, 282.9597, 283.0559, 283.1521, 283.2483, 283.3445, 283.4407, 
    283.5369, 283.6331, 283.7295, 283.8257, 283.7771, 283.6609, 283.5447, 
    283.4285, 283.3123, 283.196, 283.0796, 282.9634, 282.8472, 282.731, 
    282.6147, 282.4985, 282.3823, 282.3018, 282.2881, 282.2744, 282.2607, 
    282.2473, 282.2336, 282.22, 282.2063, 282.1926, 282.1792, 282.1655, 
    282.1519, 282.1382, 282.1245, 282.0999, 282.0754, 282.0508, 282.0264, 
    282.0017, 281.9773, 281.9526, 281.9282, 281.9036, 281.8792, 281.8547, 
    281.8301, 281.8057, 281.751, 281.6821, 281.6133, 281.5447, 281.4758, 
    281.4072, 281.3384, 281.2695, 281.2009, 281.1321, 281.0635, 280.9946, 
    280.926, 280.8665, 280.8242, 280.782, 280.7395, 280.6973, 280.655, 
    280.6128, 280.5706, 280.5283, 280.4861, 280.4438, 280.4016, 280.3591, 
    280.3176, 280.313, 280.3086, 280.304, 280.2993, 280.2949, 280.2903, 
    280.2856, 280.2812, 280.2766, 280.2722, 280.2676, 280.2629, 280.2585, 
    280.231, 280.1926, 280.1543, 280.116, 280.0776, 280.0393, 280.0012, 
    279.9629, 279.9246, 279.8862, 279.8479, 279.8096, 279.7712, 279.7349, 
    279.7017, 279.6687, 279.6355, 279.6025, 279.5693, 279.5364, 279.5032, 
    279.4702, 279.437, 279.4041, 279.3708, 279.3379, 279.3054, 279.3176, 
    279.3301, 279.3423, 279.3545, 279.3667, 279.3789, 279.3911, 279.4036, 
    279.4158, 279.428, 279.4402, 279.4524, 279.4646, 279.4573, 279.4409, 
    279.4243, 279.408, 279.3914, 279.375, 279.3584,
  277.1426, 277.1873, 277.2317, 277.2761, 277.3206, 277.365, 277.4097, 
    277.4541, 277.4985, 277.543, 277.5874, 277.6318, 277.7119, 277.8596, 
    278.0073, 278.155, 278.3027, 278.4504, 278.5981, 278.7458, 278.8936, 
    279.0413, 279.189, 279.3367, 279.4844, 279.6306, 279.6489, 279.667, 
    279.6853, 279.7034, 279.7217, 279.74, 279.7581, 279.7764, 279.7947, 
    279.8127, 279.8311, 279.8491, 279.8674, 279.895, 279.9272, 279.9592, 
    279.9915, 280.0234, 280.0557, 280.0876, 280.1199, 280.1519, 280.1841, 
    280.2161, 280.2483, 280.2803, 280.3477, 280.4819, 280.6162, 280.7505, 
    280.8848, 281.0188, 281.1531, 281.2874, 281.4216, 281.5559, 281.6902, 
    281.8245, 281.9587, 282.0918, 282.1382, 282.1846, 282.231, 282.2776, 
    282.324, 282.3704, 282.4167, 282.4631, 282.5095, 282.5559, 282.6023, 
    282.6487, 282.6951, 282.6804, 282.637, 282.5935, 282.5498, 282.5063, 
    282.4629, 282.4194, 282.3757, 282.3323, 282.2888, 282.2454, 282.2017, 
    282.1582, 282.1467, 282.1956, 282.2444, 282.2935, 282.3423, 282.3911, 
    282.4399, 282.489, 282.5378, 282.5867, 282.6355, 282.6846, 282.7334, 
    282.7815, 282.7661, 282.7505, 282.7344, 282.7178, 282.7004, 282.6829, 
    282.6646, 282.6458, 282.6265, 282.6062, 282.5857, 282.5642, 282.542, 
    282.4663, 282.3687, 282.2742, 282.1826, 282.0942, 282.0085, 281.9255, 
    281.8452, 281.7673, 281.6917, 281.6182, 281.5469, 281.4775, 281.4634, 
    281.55, 281.6365, 281.7229, 281.8093, 281.8958, 281.9824, 282.0688, 
    282.1553, 282.2417, 282.3281, 282.4148, 282.5012, 282.5876, 282.6821, 
    282.7766, 282.8711, 282.9653, 283.0598, 283.1543, 283.2485, 283.343, 
    283.4375, 283.5317, 283.6262, 283.7207, 283.8152, 283.7651, 283.6475, 
    283.5295, 283.4119, 283.2942, 283.1765, 283.0588, 282.9412, 282.8235, 
    282.7058, 282.5879, 282.4702, 282.3525, 282.2708, 282.2556, 282.2407, 
    282.2258, 282.2109, 282.1958, 282.1809, 282.166, 282.1511, 282.136, 
    282.1211, 282.1062, 282.0913, 282.0762, 282.053, 282.03, 282.0068, 
    281.9839, 281.9607, 281.9377, 281.9146, 281.8916, 281.8684, 281.8455, 
    281.8223, 281.7993, 281.7761, 281.7244, 281.6592, 281.5938, 281.5286, 
    281.4634, 281.3982, 281.333, 281.2676, 281.2024, 281.1372, 281.072, 
    281.0066, 280.9414, 280.8831, 280.8372, 280.7915, 280.7458, 280.7002, 
    280.6543, 280.6086, 280.563, 280.5171, 280.4714, 280.4258, 280.3801, 
    280.3342, 280.2893, 280.2866, 280.2842, 280.2817, 280.2791, 280.2766, 
    280.2739, 280.2715, 280.2688, 280.2664, 280.2639, 280.2612, 280.2588, 
    280.2561, 280.2324, 280.1987, 280.165, 280.1311, 280.0974, 280.0637, 
    280.03, 279.9963, 279.9626, 279.929, 279.8953, 279.8616, 279.8279, 
    279.7937, 279.7585, 279.7234, 279.6885, 279.6533, 279.6184, 279.5833, 
    279.5481, 279.5132, 279.478, 279.4429, 279.408, 279.3728, 279.3384, 
    279.3423, 279.3462, 279.3501, 279.354, 279.3579, 279.3618, 279.3657, 
    279.3696, 279.3735, 279.3774, 279.3813, 279.3853, 279.3892, 279.3848, 
    279.3765, 279.3682, 279.3599, 279.3516, 279.3433, 279.335,
  277.1624, 277.2004, 277.2385, 277.2764, 277.3145, 277.3525, 277.3906, 
    277.4287, 277.4668, 277.5049, 277.543, 277.5811, 277.6548, 277.7966, 
    277.9385, 278.0803, 278.2222, 278.3638, 278.5056, 278.6475, 278.7893, 
    278.9312, 279.073, 279.2146, 279.3564, 279.4971, 279.5317, 279.5662, 
    279.6006, 279.6353, 279.6697, 279.7043, 279.7388, 279.7732, 279.8079, 
    279.8423, 279.8767, 279.9114, 279.9458, 279.9648, 279.9768, 279.9885, 
    280.0002, 280.012, 280.0239, 280.0356, 280.0474, 280.0591, 280.071, 
    280.0828, 280.0945, 280.1062, 280.1614, 280.2991, 280.4365, 280.5742, 
    280.7117, 280.8494, 280.9868, 281.1245, 281.262, 281.3997, 281.5371, 
    281.6748, 281.8123, 281.949, 282.0156, 282.082, 282.1487, 282.2151, 
    282.2817, 282.3481, 282.4148, 282.4812, 282.5479, 282.6143, 282.6809, 
    282.7473, 282.814, 282.79, 282.7236, 282.6572, 282.5906, 282.5242, 
    282.4575, 282.3911, 282.3247, 282.2581, 282.1917, 282.125, 282.0586, 
    281.9922, 281.9753, 282.0522, 282.1294, 282.2065, 282.2834, 282.3606, 
    282.4377, 282.5146, 282.5918, 282.6689, 282.7458, 282.823, 282.9001, 
    282.9758, 282.959, 282.9409, 282.9221, 282.9026, 282.8818, 282.8601, 
    282.8372, 282.8127, 282.7871, 282.76, 282.7312, 282.7007, 282.6682, 
    282.5903, 282.4968, 282.4092, 282.3264, 282.2483, 282.1746, 282.1047, 
    282.0386, 281.9756, 281.916, 281.8591, 281.8049, 281.7532, 281.7437, 
    281.8096, 281.8755, 281.9414, 282.0073, 282.0732, 282.1392, 282.2051, 
    282.271, 282.3369, 282.4026, 282.4685, 282.5344, 282.6008, 282.6934, 
    282.7859, 282.8787, 282.9712, 283.0637, 283.1562, 283.249, 283.3416, 
    283.4341, 283.5269, 283.6194, 283.7119, 283.8044, 283.7529, 283.6338, 
    283.5146, 283.3955, 283.2764, 283.1572, 283.0378, 282.9187, 282.7996, 
    282.6804, 282.5613, 282.4421, 282.323, 282.2395, 282.2234, 282.207, 
    282.1907, 282.1746, 282.1582, 282.1418, 282.1255, 282.1094, 282.093, 
    282.0767, 282.0605, 282.0442, 282.0278, 282.0061, 281.9846, 281.9629, 
    281.9414, 281.9197, 281.8982, 281.8765, 281.855, 281.8333, 281.8118, 
    281.79, 281.7686, 281.7468, 281.6978, 281.636, 281.5745, 281.5127, 
    281.4509, 281.3892, 281.3274, 281.2656, 281.2039, 281.1421, 281.0803, 
    281.0186, 280.957, 280.8997, 280.8503, 280.8013, 280.752, 280.7029, 
    280.6536, 280.6045, 280.5552, 280.5061, 280.457, 280.4077, 280.3586, 
    280.3093, 280.261, 280.2605, 280.2598, 280.2593, 280.2588, 280.2583, 
    280.2578, 280.2571, 280.2566, 280.2561, 280.2556, 280.2549, 280.2544, 
    280.2539, 280.2339, 280.2046, 280.1755, 280.1465, 280.1174, 280.0881, 
    280.0591, 280.03, 280.0007, 279.9717, 279.9426, 279.9133, 279.8843, 
    279.8523, 279.8154, 279.7783, 279.7412, 279.7041, 279.6672, 279.6301, 
    279.593, 279.5559, 279.519, 279.4819, 279.4448, 279.4077, 279.3713, 
    279.3669, 279.3625, 279.3582, 279.3535, 279.3491, 279.3447, 279.3403, 
    279.3359, 279.3315, 279.3271, 279.3228, 279.3181, 279.3137, 279.3123, 
    279.312, 279.312, 279.3118, 279.3115, 279.3115, 279.3113,
  277.1819, 277.2134, 277.2451, 277.2769, 277.3086, 277.3403, 277.3718, 
    277.4036, 277.4353, 277.467, 277.4985, 277.5303, 277.5979, 277.7336, 
    277.8696, 278.0056, 278.1414, 278.2773, 278.4133, 278.5491, 278.6851, 
    278.821, 278.9568, 279.0928, 279.2288, 279.3638, 279.4146, 279.4653, 
    279.5161, 279.5669, 279.6177, 279.6685, 279.7192, 279.7703, 279.821, 
    279.8718, 279.9226, 279.9734, 280.0242, 280.0349, 280.0264, 280.0178, 
    280.0093, 280.0007, 279.9922, 279.9836, 279.9751, 279.9666, 279.958, 
    279.9495, 279.9409, 279.9324, 279.9753, 280.1162, 280.2571, 280.3979, 
    280.5388, 280.6797, 280.8206, 280.9614, 281.1023, 281.2432, 281.384, 
    281.5251, 281.666, 281.8062, 281.8928, 281.9795, 282.0662, 282.1528, 
    282.2395, 282.3262, 282.4128, 282.4995, 282.5862, 282.6729, 282.7595, 
    282.8462, 282.9329, 282.8999, 282.8103, 282.7209, 282.6313, 282.542, 
    282.4524, 282.3628, 282.2734, 282.1838, 282.0945, 282.0049, 281.9155, 
    281.8259, 281.804, 281.9092, 282.0144, 282.1196, 282.2249, 282.3301, 
    282.4353, 282.5405, 282.6458, 282.751, 282.8562, 282.9617, 283.0669, 
    283.1704, 283.155, 283.1384, 283.1208, 283.1018, 283.0815, 283.0596, 
    283.0359, 283.0103, 282.9824, 282.9519, 282.9187, 282.8821, 282.8416, 
    282.7588, 282.6655, 282.5811, 282.5039, 282.4336, 282.3689, 282.3096, 
    282.2544, 282.2036, 282.156, 282.1121, 282.0708, 282.032, 282.0239, 
    282.0691, 282.1145, 282.1599, 282.2053, 282.2505, 282.2959, 282.3413, 
    282.3865, 282.4319, 282.4773, 282.5225, 282.5679, 282.6138, 282.7046, 
    282.7954, 282.8862, 282.9771, 283.0676, 283.1584, 283.2493, 283.3401, 
    283.4309, 283.5217, 283.6125, 283.7031, 283.7939, 283.7407, 283.6201, 
    283.4995, 283.3789, 283.2583, 283.1377, 283.0171, 282.8965, 282.7759, 
    282.6553, 282.5347, 282.4141, 282.2935, 282.2085, 282.1909, 282.1733, 
    282.1558, 282.1382, 282.1204, 282.1028, 282.0852, 282.0676, 282.05, 
    282.0325, 282.0146, 281.9971, 281.9795, 281.9592, 281.9392, 281.9189, 
    281.8989, 281.8787, 281.8586, 281.8384, 281.8181, 281.7981, 281.7778, 
    281.7578, 281.7375, 281.7175, 281.6714, 281.613, 281.5549, 281.4966, 
    281.4385, 281.3801, 281.3218, 281.2637, 281.2053, 281.1472, 281.0889, 
    281.0308, 280.9724, 280.9163, 280.8635, 280.8108, 280.7583, 280.7056, 
    280.6528, 280.6003, 280.5476, 280.4949, 280.4424, 280.3896, 280.3372, 
    280.2844, 280.2327, 280.2341, 280.2356, 280.2371, 280.2385, 280.24, 
    280.2415, 280.2429, 280.2444, 280.2458, 280.2473, 280.2488, 280.2502, 
    280.2517, 280.2354, 280.2107, 280.1863, 280.1616, 280.1372, 280.1125, 
    280.0881, 280.0635, 280.0391, 280.0144, 279.99, 279.9653, 279.9407, 
    279.9111, 279.8721, 279.833, 279.7942, 279.7551, 279.7161, 279.677, 
    279.6379, 279.5989, 279.5598, 279.521, 279.4819, 279.4429, 279.4043, 
    279.3916, 279.3787, 279.366, 279.3533, 279.3403, 279.3276, 279.3149, 
    279.3022, 279.2893, 279.2766, 279.2639, 279.2512, 279.2383, 279.2397, 
    279.2478, 279.2556, 279.2637, 279.2717, 279.2795, 279.2876,
  277.2014, 277.2266, 277.252, 277.2771, 277.3025, 277.3279, 277.353, 
    277.3784, 277.4036, 277.429, 277.4541, 277.4795, 277.5408, 277.6709, 
    277.8008, 277.9309, 278.0608, 278.1909, 278.3208, 278.4509, 278.5808, 
    278.7109, 278.8408, 278.9709, 279.1008, 279.2302, 279.2974, 279.3645, 
    279.4314, 279.4985, 279.5657, 279.6328, 279.7, 279.7671, 279.8342, 
    279.9014, 279.9685, 280.0354, 280.1025, 280.1047, 280.0759, 280.0469, 
    280.0181, 279.9893, 279.9604, 279.9314, 279.9026, 279.8738, 279.845, 
    279.8162, 279.7871, 279.7583, 279.7891, 279.9333, 280.0776, 280.2217, 
    280.366, 280.5103, 280.6543, 280.7986, 280.9426, 281.0869, 281.2312, 
    281.3752, 281.5195, 281.6633, 281.77, 281.877, 281.9836, 282.0906, 
    282.1973, 282.304, 282.4109, 282.5176, 282.6245, 282.7312, 282.8381, 
    282.9448, 283.0518, 283.0095, 282.897, 282.7847, 282.6721, 282.5596, 
    282.4473, 282.3347, 282.2222, 282.1096, 281.9973, 281.8848, 281.7722, 
    281.6599, 281.6323, 281.7659, 281.8992, 282.0327, 282.166, 282.2996, 
    282.4329, 282.5664, 282.6997, 282.8333, 282.9666, 283.1001, 283.2334, 
    283.365, 283.3547, 283.3433, 283.3308, 283.3174, 283.3025, 283.2859, 
    283.2678, 283.2473, 283.2244, 283.1985, 283.1689, 283.1348, 283.095, 
    283.0002, 282.8965, 282.8069, 282.729, 282.6606, 282.5999, 282.5459, 
    282.4973, 282.4536, 282.4138, 282.3777, 282.3445, 282.314, 282.304, 
    282.3289, 282.3535, 282.3784, 282.4031, 282.428, 282.4526, 282.4773, 
    282.5022, 282.5269, 282.5518, 282.5764, 282.6013, 282.627, 282.7158, 
    282.8047, 282.8938, 282.9827, 283.0718, 283.1606, 283.2498, 283.3386, 
    283.4275, 283.5166, 283.6055, 283.6946, 283.7834, 283.7288, 283.6067, 
    283.4846, 283.3625, 283.2405, 283.1184, 282.9963, 282.8743, 282.752, 
    282.6299, 282.5078, 282.3857, 282.2637, 282.1775, 282.1587, 282.1396, 
    282.1206, 282.1018, 282.0828, 282.0637, 282.0449, 282.0259, 282.0068, 
    281.988, 281.969, 281.9502, 281.9312, 281.9124, 281.8938, 281.875, 
    281.8564, 281.8376, 281.8188, 281.8003, 281.7815, 281.7629, 281.7441, 
    281.7256, 281.7068, 281.688, 281.6448, 281.5901, 281.5354, 281.4807, 
    281.4258, 281.3711, 281.3164, 281.2617, 281.2068, 281.1521, 281.0974, 
    281.0427, 280.988, 280.9326, 280.8767, 280.8206, 280.7644, 280.7083, 
    280.6521, 280.5962, 280.54, 280.4839, 280.4277, 280.3716, 280.3157, 
    280.2595, 280.2043, 280.2078, 280.2112, 280.2146, 280.2183, 280.2217, 
    280.2251, 280.2285, 280.2319, 280.2354, 280.239, 280.2424, 280.2458, 
    280.2493, 280.2368, 280.2168, 280.1968, 280.177, 280.157, 280.137, 
    280.1169, 280.0972, 280.0771, 280.0571, 280.0371, 280.0173, 279.9973, 
    279.97, 279.929, 279.8879, 279.8469, 279.8059, 279.7649, 279.7239, 
    279.6829, 279.6418, 279.6008, 279.5598, 279.5188, 279.4778, 279.4373, 
    279.416, 279.395, 279.3738, 279.3528, 279.3318, 279.3105, 279.2896, 
    279.2683, 279.2473, 279.2261, 279.2051, 279.1841, 279.1628, 279.1672, 
    279.1833, 279.1995, 279.2156, 279.2317, 279.2478, 279.2639,
  277.2209, 277.2397, 277.2588, 277.2776, 277.2964, 277.3154, 277.3342, 
    277.353, 277.3721, 277.3909, 277.4097, 277.4287, 277.4836, 277.6079, 
    277.7319, 277.856, 277.9802, 278.1042, 278.2283, 278.3525, 278.4766, 
    278.6006, 278.7249, 278.8489, 278.9729, 279.0967, 279.1802, 279.2634, 
    279.3469, 279.4304, 279.5137, 279.5972, 279.6807, 279.7639, 279.8474, 
    279.9309, 280.0142, 280.0977, 280.1809, 280.1746, 280.1252, 280.0762, 
    280.0271, 279.9778, 279.9287, 279.8794, 279.8303, 279.781, 279.7319, 
    279.6826, 279.6335, 279.5842, 279.603, 279.7505, 279.8979, 280.0457, 
    280.1931, 280.3406, 280.488, 280.6355, 280.7832, 280.9307, 281.0781, 
    281.2256, 281.373, 281.5205, 281.6472, 281.7742, 281.9011, 282.0281, 
    282.155, 282.282, 282.4089, 282.5359, 282.6628, 282.7898, 282.9167, 
    283.0437, 283.1704, 283.1194, 282.9839, 282.8484, 282.7129, 282.5774, 
    282.4419, 282.3064, 282.1709, 282.0356, 281.9001, 281.7646, 281.6292, 
    281.4937, 281.4609, 281.6226, 281.7842, 281.9458, 282.1074, 282.269, 
    282.4307, 282.5923, 282.7539, 282.9155, 283.0769, 283.2385, 283.4001, 
    283.5598, 283.5579, 283.5559, 283.5537, 283.5513, 283.5483, 283.5452, 
    283.5415, 283.5374, 283.5325, 283.5266, 283.5195, 283.5107, 283.4998, 
    283.376, 283.2327, 283.1177, 283.0237, 282.9453, 282.8789, 282.8218, 
    282.7725, 282.7292, 282.6909, 282.657, 282.6267, 282.5994, 282.5842, 
    282.5884, 282.5925, 282.5969, 282.6011, 282.6052, 282.6094, 282.6135, 
    282.6177, 282.6221, 282.6262, 282.6304, 282.6345, 282.6399, 282.7271, 
    282.8142, 282.9014, 282.9885, 283.0757, 283.1628, 283.25, 283.3372, 
    283.4243, 283.5115, 283.5986, 283.6858, 283.7729, 283.7166, 283.593, 
    283.4695, 283.3459, 283.2224, 283.0989, 282.9753, 282.8518, 282.7283, 
    282.6047, 282.4812, 282.3577, 282.2341, 282.1465, 282.1262, 282.106, 
    282.0857, 282.0654, 282.0452, 282.0249, 282.0044, 281.9841, 281.9639, 
    281.9436, 281.9233, 281.9031, 281.8828, 281.8655, 281.8484, 281.8311, 
    281.814, 281.7966, 281.7793, 281.7622, 281.7449, 281.7278, 281.7104, 
    281.6931, 281.676, 281.6587, 281.6184, 281.5671, 281.5159, 281.4646, 
    281.4133, 281.3621, 281.3108, 281.2595, 281.2085, 281.1572, 281.106, 
    281.0547, 281.0034, 280.9492, 280.8896, 280.8301, 280.7705, 280.7109, 
    280.6514, 280.5918, 280.5325, 280.4729, 280.4133, 280.3538, 280.2942, 
    280.2346, 280.176, 280.1814, 280.187, 280.1924, 280.1978, 280.2034, 
    280.2087, 280.2141, 280.2197, 280.2251, 280.2307, 280.2361, 280.2415, 
    280.2471, 280.2383, 280.2229, 280.2075, 280.1921, 280.1768, 280.1614, 
    280.146, 280.1306, 280.1152, 280.0999, 280.0845, 280.0691, 280.0537, 
    280.0288, 279.9858, 279.9429, 279.8997, 279.8567, 279.8137, 279.7708, 
    279.7278, 279.6848, 279.6418, 279.5989, 279.5559, 279.5129, 279.4702, 
    279.4407, 279.4111, 279.3818, 279.3523, 279.323, 279.2935, 279.2642, 
    279.2346, 279.2051, 279.1758, 279.1462, 279.1169, 279.0874, 279.0947, 
    279.1189, 279.1433, 279.1675, 279.1919, 279.2161, 279.2405,
  277.2405, 277.2529, 277.2654, 277.2778, 277.2905, 277.303, 277.3154, 
    277.3279, 277.3403, 277.3528, 277.3652, 277.3779, 277.4268, 277.5449, 
    277.6631, 277.7812, 277.8994, 278.0178, 278.136, 278.2542, 278.3723, 
    278.4905, 278.6089, 278.7271, 278.8452, 278.9631, 279.063, 279.1626, 
    279.2622, 279.3621, 279.4617, 279.5615, 279.6611, 279.761, 279.8606, 
    279.9602, 280.0601, 280.1597, 280.2595, 280.2444, 280.1748, 280.1055, 
    280.0359, 279.9663, 279.897, 279.8274, 279.7578, 279.6885, 279.6189, 
    279.5493, 279.48, 279.4104, 279.417, 279.5676, 279.7185, 279.8694, 
    280.0203, 280.1709, 280.3218, 280.4727, 280.6235, 280.7742, 280.925, 
    281.0759, 281.2268, 281.3774, 281.5247, 281.6716, 281.8188, 281.9658, 
    282.1128, 282.26, 282.407, 282.554, 282.7012, 282.8481, 282.9954, 
    283.1423, 283.2893, 283.229, 283.0706, 282.9121, 282.7537, 282.5952, 
    282.4368, 282.2783, 282.1199, 281.9614, 281.803, 281.6445, 281.4861, 
    281.3276, 281.2896, 281.4792, 281.6692, 281.8589, 282.0486, 282.2385, 
    282.4282, 282.6179, 282.8079, 282.9976, 283.1873, 283.3772, 283.5669, 
    283.7544, 283.7649, 283.7769, 283.7903, 283.8059, 284.5349, 284.5923, 
    284.6389, 284.6775, 284.7097, 284.7373, 284.7612, 284.7817, 284.8, 
    284.0405, 283.7666, 283.5718, 283.4258, 283.3125, 283.2222, 283.1482, 
    283.0867, 283.0344, 282.99, 282.9514, 282.9175, 282.8877, 282.8645, 
    282.8481, 282.8318, 282.8154, 282.7988, 282.7825, 282.7661, 282.7498, 
    282.7334, 282.717, 282.7007, 282.6843, 282.668, 282.6528, 282.7383, 
    282.8237, 282.9089, 282.9944, 283.0796, 283.165, 283.2502, 283.3357, 
    283.4211, 283.5063, 283.5918, 283.677, 283.7625, 283.7046, 283.5796, 
    283.4546, 283.3296, 283.2046, 283.0796, 282.9546, 282.8296, 282.7046, 
    282.5796, 282.4546, 282.3296, 282.2046, 282.1155, 282.0938, 282.0723, 
    282.0505, 282.0291, 282.0073, 281.9858, 281.9641, 281.9424, 281.9209, 
    281.8992, 281.8777, 281.856, 281.8345, 281.8186, 281.803, 281.7871, 
    281.7712, 281.7556, 281.7397, 281.7241, 281.7083, 281.6924, 281.6768, 
    281.6609, 281.6453, 281.6294, 281.5918, 281.5439, 281.4963, 281.4485, 
    281.4009, 281.353, 281.3054, 281.2576, 281.21, 281.1621, 281.1145, 
    281.0667, 281.019, 280.9658, 280.9028, 280.8398, 280.7769, 280.7139, 
    280.6509, 280.5876, 280.5247, 280.4617, 280.3987, 280.3357, 280.2727, 
    280.2097, 280.1477, 280.1553, 280.1626, 280.1702, 280.1775, 280.1851, 
    280.1924, 280.2, 280.2073, 280.2148, 280.2224, 280.2297, 280.2373, 
    280.2446, 280.2397, 280.229, 280.218, 280.2073, 280.1965, 280.1858, 
    280.175, 280.1641, 280.1533, 280.1426, 280.1318, 280.1211, 280.1104, 
    280.0874, 280.0425, 279.9976, 279.9526, 279.9077, 279.8625, 279.8176, 
    279.7727, 279.7278, 279.6829, 279.6379, 279.5928, 279.5479, 279.5029, 
    279.4653, 279.4275, 279.3896, 279.3521, 279.3142, 279.2764, 279.2385, 
    279.2009, 279.1631, 279.1252, 279.0876, 279.0498, 279.012, 279.0222, 
    279.0547, 279.0872, 279.1194, 279.1519, 279.1843, 279.2168,
  277.3057, 277.3162, 277.3267, 277.3372, 277.3477, 277.3584, 277.3689, 
    277.3794, 277.3899, 277.4004, 277.4109, 277.4216, 277.468, 277.5828, 
    277.6975, 277.8125, 277.9272, 278.0422, 278.157, 278.2717, 278.3867, 
    278.5015, 278.6165, 278.7312, 278.8459, 278.9609, 279.0735, 279.1863, 
    279.2991, 279.4116, 279.5244, 279.6372, 279.75, 279.8625, 279.9753, 
    280.0881, 280.2007, 280.3135, 280.4263, 280.4128, 280.3396, 280.2661, 
    280.1929, 280.1196, 280.0461, 279.9729, 279.8997, 279.8264, 279.7529, 
    279.6797, 279.6064, 279.5332, 279.5352, 279.6804, 279.8259, 279.9712, 
    280.1165, 280.2617, 280.407, 280.5522, 280.6975, 280.8428, 280.9883, 
    281.1335, 281.2788, 281.4243, 281.5928, 281.761, 281.9292, 282.0977, 
    282.2659, 282.4343, 282.6025, 282.7708, 282.9392, 283.1074, 283.2759, 
    283.4441, 283.6123, 283.5503, 283.3792, 283.2083, 283.0371, 282.8662, 
    282.6951, 282.5239, 282.353, 282.1819, 282.011, 281.8398, 281.6687, 
    281.4978, 281.449, 281.6313, 281.8135, 281.9958, 282.178, 282.3604, 
    282.5427, 282.7249, 282.9072, 283.0894, 283.2717, 283.4541, 283.6362, 
    283.8164, 283.8306, 283.8469, 283.8655, 283.887, 284.4854, 284.533, 
    284.5713, 284.603, 284.6296, 284.6521, 284.6714, 284.6882, 284.7031, 
    284.3137, 283.9287, 283.6719, 283.4883, 283.3503, 283.2432, 283.1572, 
    283.0872, 283.0286, 282.979, 282.9365, 282.8997, 282.8674, 282.8442, 
    282.8318, 282.8196, 282.8071, 282.7947, 282.7825, 282.77, 282.7576, 
    282.7454, 282.7329, 282.7205, 282.7083, 282.6958, 282.6848, 282.7625, 
    282.8401, 282.9177, 282.9954, 283.073, 283.1506, 283.2283, 283.3062, 
    283.3838, 283.4614, 283.5391, 283.6167, 283.6943, 283.6355, 283.5125, 
    283.3896, 283.2668, 283.1438, 283.021, 282.8979, 282.7751, 282.6523, 
    282.5293, 282.4065, 282.2837, 282.1606, 282.0718, 282.0469, 282.0217, 
    281.9968, 281.9717, 281.9468, 281.9216, 281.8965, 281.8716, 281.8464, 
    281.8215, 281.7964, 281.7715, 281.7466, 281.7332, 281.7197, 281.7065, 
    281.6931, 281.6797, 281.6665, 281.6531, 281.6396, 281.6265, 281.613, 
    281.5996, 281.5864, 281.573, 281.5391, 281.4954, 281.4519, 281.4084, 
    281.3647, 281.3213, 281.2776, 281.2341, 281.1907, 281.147, 281.1035, 
    281.0598, 281.0164, 280.9666, 280.9048, 280.8433, 280.7817, 280.72, 
    280.6584, 280.5969, 280.5352, 280.4736, 280.4121, 280.3503, 280.2888, 
    280.2273, 280.1667, 280.176, 280.1853, 280.1946, 280.2039, 280.2131, 
    280.2224, 280.2317, 280.2407, 280.25, 280.2593, 280.2686, 280.2778, 
    280.2871, 280.2837, 280.2742, 280.2646, 280.2551, 280.2456, 280.2361, 
    280.2266, 280.2173, 280.2078, 280.1982, 280.1887, 280.1792, 280.1697, 
    280.1477, 280.1028, 280.0576, 280.0125, 279.9673, 279.9221, 279.877, 
    279.8318, 279.7869, 279.7417, 279.6965, 279.6514, 279.6062, 279.5613, 
    279.5195, 279.4778, 279.436, 279.3943, 279.3525, 279.3108, 279.269, 
    279.2273, 279.1855, 279.1438, 279.1021, 279.0603, 279.0186, 279.0225, 
    279.0476, 279.0728, 279.0977, 279.1228, 279.1477, 279.1729,
  277.3977, 277.4089, 277.4202, 277.4314, 277.4426, 277.4539, 277.4651, 
    277.4763, 277.4875, 277.4988, 277.51, 277.5212, 277.5674, 277.6804, 
    277.7932, 277.9062, 278.0193, 278.1321, 278.2451, 278.3582, 278.4709, 
    278.584, 278.697, 278.8101, 278.9229, 279.0359, 279.1597, 279.2834, 
    279.4075, 279.5312, 279.655, 279.7788, 279.9026, 280.0264, 280.1501, 
    280.2739, 280.3977, 280.5215, 280.6453, 280.6394, 280.572, 280.5046, 
    280.4375, 280.3701, 280.3027, 280.2354, 280.168, 280.1006, 280.0332, 
    279.9661, 279.8987, 279.8313, 279.8335, 279.968, 280.1028, 280.2373, 
    280.3718, 280.5063, 280.6409, 280.7754, 280.9099, 281.0444, 281.179, 
    281.3135, 281.448, 281.5833, 281.7734, 281.9636, 282.1541, 282.3442, 
    282.5344, 282.7246, 282.9148, 283.105, 283.2952, 283.4854, 283.6758, 
    283.866, 284.0562, 283.9966, 283.8191, 283.6416, 283.4641, 283.2866, 
    283.1091, 282.9316, 282.7542, 282.5767, 282.3994, 282.2219, 282.0444, 
    281.8669, 281.804, 281.9575, 282.1113, 282.2649, 282.4187, 282.5723, 
    282.7261, 282.8796, 283.0334, 283.187, 283.3408, 283.4944, 283.6482, 
    283.8, 283.8113, 283.8242, 283.8389, 283.856, 284.332, 284.3699, 
    284.4006, 284.4258, 284.4468, 284.4646, 284.4802, 284.4937, 284.5054, 
    284.114, 283.7278, 283.47, 283.2859, 283.1477, 283.04, 282.9541, 
    282.8835, 282.8247, 282.7751, 282.7324, 282.6956, 282.6633, 282.6465, 
    282.6526, 282.6587, 282.665, 282.6711, 282.6772, 282.6836, 282.6897, 
    282.6958, 282.7021, 282.7083, 282.7144, 282.7207, 282.7275, 282.7942, 
    282.8606, 282.9272, 282.9937, 283.0603, 283.1267, 283.1934, 283.2598, 
    283.3262, 283.3928, 283.4592, 283.5259, 283.5923, 283.5327, 283.4141, 
    283.2954, 283.1768, 283.0579, 282.9392, 282.8206, 282.7019, 282.5833, 
    282.4646, 282.3459, 282.2273, 282.1084, 282.0208, 281.9912, 281.9614, 
    281.9316, 281.9021, 281.8723, 281.8425, 281.813, 281.7832, 281.7537, 
    281.7239, 281.6941, 281.6646, 281.635, 281.6248, 281.6145, 281.604, 
    281.5938, 281.5835, 281.573, 281.5627, 281.5522, 281.542, 281.5317, 
    281.5212, 281.511, 281.5005, 281.4707, 281.4319, 281.3928, 281.3538, 
    281.3149, 281.2759, 281.2368, 281.198, 281.1589, 281.1201, 281.0811, 
    281.042, 281.0032, 280.9578, 280.9004, 280.843, 280.7859, 280.7285, 
    280.6711, 280.6138, 280.5564, 280.4993, 280.4419, 280.3845, 280.3271, 
    280.27, 280.2136, 280.2246, 280.2356, 280.2466, 280.2576, 280.2686, 
    280.2795, 280.2903, 280.3013, 280.3123, 280.3232, 280.3342, 280.3452, 
    280.3562, 280.3525, 280.3425, 280.3323, 280.3223, 280.312, 280.302, 
    280.2917, 280.2817, 280.2715, 280.2615, 280.2512, 280.2412, 280.231, 
    280.209, 280.1648, 280.1206, 280.0764, 280.0322, 279.9878, 279.9436, 
    279.8994, 279.8552, 279.811, 279.7668, 279.7227, 279.6785, 279.6343, 
    279.5911, 279.5481, 279.5049, 279.4619, 279.4187, 279.3755, 279.3325, 
    279.2893, 279.2463, 279.2031, 279.1599, 279.1169, 279.0737, 279.0659, 
    279.0745, 279.083, 279.0913, 279.0999, 279.1084, 279.1167,
  277.4897, 277.5015, 277.5134, 277.5254, 277.5374, 277.5493, 277.561, 
    277.573, 277.585, 277.5969, 277.6089, 277.6206, 277.6667, 277.7778, 
    277.8889, 278, 278.1111, 278.2222, 278.3333, 278.4443, 278.5554, 
    278.6665, 278.7776, 278.8887, 278.9998, 279.1111, 279.2461, 279.3809, 
    279.5156, 279.6506, 279.7854, 279.9202, 280.0552, 280.1899, 280.325, 
    280.4597, 280.5945, 280.7295, 280.8643, 280.866, 280.8047, 280.7432, 
    280.6819, 280.6206, 280.5591, 280.4978, 280.4363, 280.375, 280.3135, 
    280.2522, 280.1909, 280.1294, 280.1318, 280.2556, 280.3794, 280.5032, 
    280.6272, 280.751, 280.8748, 280.9985, 281.1223, 281.2461, 281.3699, 
    281.4937, 281.6174, 281.7422, 281.9543, 282.1665, 282.3787, 282.5908, 
    282.8027, 283.0149, 283.2271, 283.4392, 283.6514, 283.8635, 284.0757, 
    284.2876, 284.4998, 284.4431, 284.259, 284.0752, 283.8914, 283.7073, 
    283.5234, 283.3394, 283.1555, 282.9717, 282.7876, 282.6038, 282.4199, 
    282.2358, 282.1589, 282.2839, 282.4092, 282.5342, 282.6592, 282.7844, 
    282.9094, 283.0344, 283.1597, 283.2847, 283.4097, 283.5349, 283.6599, 
    283.7834, 283.792, 283.8015, 283.8125, 283.8252, 284.179, 284.207, 
    284.2297, 284.2483, 284.2642, 284.2773, 284.2888, 284.2988, 284.3076, 
    283.9141, 283.5269, 283.2683, 283.0835, 282.9448, 282.8369, 282.7507, 
    282.6799, 282.6211, 282.5713, 282.5286, 282.4915, 282.459, 282.4487, 
    282.4734, 282.498, 282.5227, 282.5476, 282.5723, 282.5969, 282.6218, 
    282.6465, 282.6711, 282.696, 282.7207, 282.7454, 282.7705, 282.8259, 
    282.8813, 282.9368, 282.9919, 283.0474, 283.1028, 283.1582, 283.2134, 
    283.2688, 283.3242, 283.3796, 283.4348, 283.4902, 283.4299, 283.3154, 
    283.2009, 283.0867, 282.9722, 282.8577, 282.7432, 282.6287, 282.5142, 
    282.3997, 282.2852, 282.1707, 282.0564, 281.9697, 281.9353, 281.9011, 
    281.8667, 281.8323, 281.7981, 281.7637, 281.7292, 281.6951, 281.6606, 
    281.6262, 281.592, 281.5576, 281.5237, 281.5164, 281.509, 281.5017, 
    281.4944, 281.4871, 281.4797, 281.4724, 281.4648, 281.4575, 281.4502, 
    281.4429, 281.4355, 281.4282, 281.4023, 281.3682, 281.3337, 281.2993, 
    281.2649, 281.2305, 281.196, 281.1619, 281.1274, 281.093, 281.0586, 
    281.0242, 280.9897, 280.949, 280.896, 280.843, 280.7898, 280.7368, 
    280.6838, 280.6309, 280.5779, 280.5247, 280.4717, 280.4187, 280.3657, 
    280.3127, 280.2607, 280.2734, 280.2859, 280.2986, 280.3113, 280.324, 
    280.3364, 280.3491, 280.3618, 280.3745, 280.3872, 280.3997, 280.4124, 
    280.425, 280.4216, 280.4109, 280.4001, 280.3894, 280.3787, 280.3677, 
    280.3569, 280.3462, 280.3354, 280.3247, 280.314, 280.303, 280.2922, 
    280.2703, 280.2268, 280.1836, 280.1404, 280.0969, 280.0537, 280.0105, 
    279.967, 279.9238, 279.8806, 279.8372, 279.7939, 279.7507, 279.7073, 
    279.6628, 279.6184, 279.5737, 279.5293, 279.4849, 279.4404, 279.396, 
    279.3513, 279.3069, 279.2625, 279.218, 279.1736, 279.1289, 279.1094, 
    279.1013, 279.0933, 279.085, 279.0769, 279.0688, 279.0608,
  277.5815, 277.5942, 277.6069, 277.6194, 277.6321, 277.6448, 277.6572, 
    277.6699, 277.6824, 277.6951, 277.7078, 277.7202, 277.7661, 277.8752, 
    277.9846, 278.0938, 278.2029, 278.3123, 278.4214, 278.5305, 278.6399, 
    278.749, 278.8582, 278.9675, 279.0767, 279.1863, 279.3323, 279.478, 
    279.624, 279.77, 279.916, 280.0618, 280.2078, 280.3538, 280.4995, 
    280.6455, 280.7915, 280.9373, 281.0833, 281.0928, 281.0374, 280.9819, 
    280.9265, 280.8711, 280.8157, 280.7603, 280.7048, 280.6492, 280.5938, 
    280.5383, 280.4829, 280.4275, 280.4302, 280.5432, 280.6562, 280.7693, 
    280.8823, 280.9954, 281.1084, 281.2214, 281.3345, 281.4475, 281.5605, 
    281.6736, 281.7866, 281.9011, 282.1353, 282.3691, 282.6033, 282.8372, 
    283.0713, 283.3054, 283.5393, 283.7734, 284.0073, 284.2415, 284.4753, 
    284.7095, 284.9436, 284.8894, 284.699, 284.5085, 284.3184, 284.1279, 
    283.9375, 283.7471, 283.5569, 283.3665, 283.176, 282.9858, 282.7954, 
    282.605, 282.5139, 282.6104, 282.7068, 282.8035, 282.8999, 282.9963, 
    283.0928, 283.1892, 283.2859, 283.3823, 283.4788, 283.5752, 283.6719, 
    283.7671, 283.7727, 283.7788, 283.7861, 283.7944, 284.0256, 284.0439, 
    284.0588, 284.071, 284.0813, 284.0901, 284.0974, 284.104, 284.1096, 
    283.7141, 283.3257, 283.0664, 282.8811, 282.7422, 282.634, 282.5474, 
    282.4766, 282.4175, 282.3674, 282.3245, 282.2874, 282.2549, 282.2507, 
    282.2942, 282.3374, 282.3806, 282.4238, 282.4673, 282.5105, 282.5537, 
    282.5972, 282.6404, 282.6836, 282.7268, 282.7703, 282.8135, 282.8577, 
    282.9019, 282.946, 282.9902, 283.0344, 283.0789, 283.123, 283.1672, 
    283.2114, 283.2556, 283.2998, 283.344, 283.3882, 283.3271, 283.217, 
    283.1067, 282.9963, 282.8862, 282.7759, 282.6658, 282.5554, 282.4451, 
    282.335, 282.2246, 282.1143, 282.0042, 281.9187, 281.8796, 281.8406, 
    281.8018, 281.7627, 281.7236, 281.6848, 281.6458, 281.6067, 281.5679, 
    281.5288, 281.4897, 281.4509, 281.4124, 281.408, 281.4036, 281.3994, 
    281.395, 281.3906, 281.3862, 281.3818, 281.3777, 281.3733, 281.3689, 
    281.3645, 281.3601, 281.356, 281.3342, 281.3044, 281.2747, 281.2449, 
    281.2148, 281.1851, 281.1553, 281.1255, 281.0957, 281.0659, 281.0361, 
    281.0063, 280.9766, 280.9402, 280.8914, 280.8428, 280.7939, 280.7454, 
    280.6965, 280.6477, 280.5991, 280.5503, 280.5017, 280.4529, 280.4041, 
    280.3555, 280.3076, 280.322, 280.3364, 280.3506, 280.365, 280.3794, 
    280.3936, 280.408, 280.4224, 280.4368, 280.4509, 280.4653, 280.4797, 
    280.4939, 280.4907, 280.4792, 280.4678, 280.4565, 280.4451, 280.4336, 
    280.4221, 280.4106, 280.3992, 280.3879, 280.3765, 280.365, 280.3535, 
    280.3313, 280.2891, 280.2466, 280.2041, 280.1619, 280.1194, 280.0771, 
    280.0347, 279.9924, 279.95, 279.9075, 279.8652, 279.8228, 279.7803, 
    279.7346, 279.6887, 279.6428, 279.5969, 279.551, 279.5051, 279.4592, 
    279.4136, 279.3677, 279.3218, 279.2759, 279.23, 279.1841, 279.1528, 
    279.1282, 279.1035, 279.0789, 279.0542, 279.0295, 279.0049,
  277.6736, 277.687, 277.7002, 277.7136, 277.7268, 277.7402, 277.7534, 
    277.7666, 277.78, 277.7932, 277.8066, 277.8198, 277.8655, 277.9729, 
    278.0801, 278.1875, 278.2949, 278.4021, 278.5095, 278.6169, 278.7241, 
    278.8315, 278.939, 279.0461, 279.1536, 279.2615, 279.4185, 279.5754, 
    279.7324, 279.8894, 280.0464, 280.2034, 280.3604, 280.5173, 280.6743, 
    280.8313, 280.9883, 281.1453, 281.3022, 281.3193, 281.2698, 281.2205, 
    281.1709, 281.1213, 281.072, 281.0225, 280.9731, 280.9236, 280.874, 
    280.8247, 280.7751, 280.7258, 280.7288, 280.8308, 280.9331, 281.0354, 
    281.1377, 281.24, 281.3423, 281.4446, 281.5469, 281.6492, 281.7515, 
    281.8538, 281.9561, 282.0601, 282.3159, 282.572, 282.8279, 283.0837, 
    283.3398, 283.5957, 283.8516, 284.1077, 284.3635, 284.6194, 284.8752, 
    285.1313, 285.3872, 285.3357, 285.1389, 284.9421, 284.7454, 284.5486, 
    284.3518, 284.1548, 283.958, 283.7612, 283.5645, 283.3677, 283.1709, 
    282.9741, 282.8689, 282.9368, 283.0046, 283.0725, 283.1404, 283.2083, 
    283.2761, 283.3442, 283.4121, 283.48, 283.5479, 283.6157, 283.6836, 
    283.7507, 283.7532, 283.7561, 283.7595, 283.7634, 283.8723, 283.8811, 
    283.8879, 283.8938, 283.8984, 283.9026, 283.9062, 283.9092, 283.9119, 
    283.5144, 283.1248, 282.8647, 282.679, 282.5393, 282.4309, 282.344, 
    282.2729, 282.2136, 282.1636, 282.1206, 282.0833, 282.0508, 282.053, 
    282.1147, 282.1768, 282.2385, 282.3003, 282.3621, 282.4241, 282.4858, 
    282.5476, 282.6094, 282.6714, 282.7332, 282.7949, 282.8564, 282.8894, 
    282.9226, 282.9556, 282.9888, 283.0217, 283.0547, 283.0879, 283.1208, 
    283.1541, 283.187, 283.22, 283.2532, 283.2861, 283.2246, 283.1184, 
    283.0125, 282.9062, 282.8003, 282.6943, 282.5881, 282.4822, 282.376, 
    282.27, 282.1641, 282.0579, 281.9519, 281.8674, 281.824, 281.7803, 
    281.7366, 281.6931, 281.6494, 281.6057, 281.562, 281.5186, 281.4749, 
    281.4312, 281.3877, 281.344, 281.301, 281.2996, 281.2983, 281.2969, 
    281.2957, 281.2942, 281.293, 281.2915, 281.2903, 281.2888, 281.2876, 
    281.2861, 281.2849, 281.2834, 281.2659, 281.2407, 281.2153, 281.1902, 
    281.165, 281.1399, 281.1145, 281.0894, 281.0642, 281.0391, 281.0137, 
    280.9885, 280.9634, 280.9314, 280.887, 280.8425, 280.7981, 280.7537, 
    280.7092, 280.6648, 280.6204, 280.5759, 280.5315, 280.4871, 280.4426, 
    280.3982, 280.3547, 280.3706, 280.3867, 280.4028, 280.4187, 280.4348, 
    280.4507, 280.4668, 280.4829, 280.4988, 280.5149, 280.5308, 280.5469, 
    280.563, 280.5598, 280.5476, 280.5356, 280.5234, 280.5115, 280.4993, 
    280.4873, 280.4753, 280.4631, 280.4512, 280.439, 280.427, 280.4148, 
    280.3926, 280.3511, 280.3096, 280.2681, 280.2266, 280.1853, 280.1438, 
    280.1023, 280.0608, 280.0193, 279.9778, 279.9365, 279.895, 279.8535, 
    279.8062, 279.759, 279.7117, 279.6646, 279.6172, 279.5701, 279.5227, 
    279.4756, 279.4282, 279.3811, 279.3337, 279.2866, 279.2393, 279.1963, 
    279.155, 279.1138, 279.0725, 279.0312, 278.99, 278.9487,
  277.7656, 277.7798, 277.7937, 277.8076, 277.8215, 277.8357, 277.8496, 
    277.8635, 277.8774, 277.8916, 277.9055, 277.9194, 277.9648, 278.0703, 
    278.1758, 278.2812, 278.3867, 278.4922, 278.5977, 278.7031, 278.8086, 
    278.9141, 279.0195, 279.125, 279.2305, 279.3367, 279.5046, 279.6726, 
    279.8408, 280.0088, 280.1768, 280.345, 280.5129, 280.6812, 280.8491, 
    281.0171, 281.1853, 281.3533, 281.5212, 281.5459, 281.5024, 281.459, 
    281.4155, 281.3718, 281.3284, 281.2849, 281.2415, 281.198, 281.1543, 
    281.1108, 281.0674, 281.0239, 281.0271, 281.1184, 281.21, 281.3015, 
    281.3931, 281.4846, 281.5762, 281.6677, 281.7593, 281.8506, 281.9421, 
    282.0337, 282.1252, 282.219, 282.4968, 282.7747, 283.0525, 283.3303, 
    283.6082, 283.886, 284.1638, 284.4417, 284.7195, 284.9973, 285.2751, 
    285.553, 285.8308, 285.782, 285.5789, 285.3755, 285.1724, 284.969, 
    284.7659, 284.5625, 284.3594, 284.1562, 283.9529, 283.7498, 283.5464, 
    283.3433, 283.2239, 283.2632, 283.3025, 283.3418, 283.3811, 283.4204, 
    283.4597, 283.499, 283.5383, 283.5776, 283.6169, 283.6562, 283.6956, 
    283.7341, 283.7339, 283.7336, 283.7332, 283.7327, 283.719, 283.718, 
    283.717, 283.7163, 283.7158, 283.7153, 283.7148, 283.7146, 283.7141, 
    283.3145, 282.9238, 282.6628, 282.4766, 282.3367, 282.2278, 282.1406, 
    282.0693, 282.01, 281.9597, 281.9165, 281.8792, 281.8464, 281.8552, 
    281.9355, 282.0159, 282.0964, 282.1768, 282.2571, 282.3374, 282.418, 
    282.4983, 282.5786, 282.6589, 282.7395, 282.8198, 282.8994, 282.9211, 
    282.9431, 282.9651, 282.9871, 283.0088, 283.0308, 283.0527, 283.0747, 
    283.0964, 283.1184, 283.1404, 283.1624, 283.1841, 283.1218, 283.02, 
    282.9182, 282.8162, 282.7144, 282.6125, 282.5107, 282.4089, 282.3071, 
    282.2051, 282.1033, 282.0015, 281.8997, 281.8164, 281.7681, 281.72, 
    281.6716, 281.6233, 281.575, 281.5269, 281.4785, 281.4302, 281.3818, 
    281.3337, 281.2854, 281.2371, 281.1895, 281.1912, 281.1929, 281.1946, 
    281.1963, 281.1978, 281.1995, 281.2012, 281.2029, 281.2046, 281.2061, 
    281.2078, 281.2095, 281.2112, 281.1975, 281.177, 281.1562, 281.1357, 
    281.115, 281.0945, 281.0737, 281.0532, 281.0325, 281.012, 280.9912, 
    280.9707, 280.95, 280.9226, 280.8826, 280.8423, 280.8022, 280.762, 
    280.7219, 280.6816, 280.6416, 280.6016, 280.5613, 280.5212, 280.481, 
    280.4409, 280.4016, 280.4194, 280.437, 280.4548, 280.4724, 280.4902, 
    280.5078, 280.5256, 280.5432, 280.561, 280.5786, 280.5964, 280.614, 
    280.6318, 280.6287, 280.616, 280.6033, 280.5906, 280.5779, 280.5652, 
    280.5525, 280.5398, 280.5271, 280.5144, 280.5015, 280.4888, 280.4761, 
    280.4536, 280.4131, 280.3726, 280.332, 280.2915, 280.251, 280.2104, 
    280.1699, 280.1294, 280.0889, 280.0483, 280.0078, 279.9673, 279.9265, 
    279.8779, 279.8293, 279.7808, 279.7319, 279.6833, 279.6348, 279.5862, 
    279.5376, 279.489, 279.4404, 279.3918, 279.343, 279.2944, 279.2395, 
    279.1819, 279.124, 279.0662, 279.0083, 278.9507, 278.8928,
  277.8577, 277.8723, 277.887, 277.9016, 277.9165, 277.9312, 277.9458, 
    277.9604, 277.9751, 277.9897, 278.0044, 278.019, 278.0642, 278.168, 
    278.2715, 278.375, 278.4788, 278.5823, 278.6858, 278.7893, 278.8931, 
    278.9966, 279.1001, 279.2039, 279.3074, 279.4119, 279.5908, 279.77, 
    279.9492, 280.1282, 280.3074, 280.4866, 280.6655, 280.8447, 281.0239, 
    281.2029, 281.3821, 281.5613, 281.7402, 281.7725, 281.7351, 281.6975, 
    281.6599, 281.6223, 281.585, 281.5474, 281.5098, 281.4722, 281.4348, 
    281.3972, 281.3596, 281.322, 281.3254, 281.406, 281.4868, 281.5676, 
    281.6484, 281.7292, 281.8101, 281.8906, 281.9714, 282.0522, 282.1331, 
    282.2139, 282.2947, 282.3779, 282.6777, 282.9775, 283.2771, 283.5769, 
    283.8767, 284.1765, 284.4761, 284.7759, 285.0757, 285.3755, 285.675, 
    285.9749, 286.2747, 286.2285, 286.0188, 285.8091, 285.5994, 285.3896, 
    285.1799, 284.9705, 284.7607, 284.551, 284.3413, 284.1316, 283.9219, 
    283.7122, 283.5789, 283.5896, 283.6001, 283.6108, 283.6216, 283.6323, 
    283.6431, 283.6538, 283.6646, 283.675, 283.6858, 283.6965, 283.7073, 
    283.7178, 283.7146, 283.7109, 283.7065, 283.7017, 283.5659, 283.5549, 
    283.5464, 283.5391, 283.533, 283.5278, 283.5234, 283.5198, 283.5164, 
    283.1145, 282.7227, 282.4612, 282.2742, 282.1338, 282.0247, 281.9373, 
    281.866, 281.8064, 281.7559, 281.7126, 281.675, 281.6423, 281.6575, 
    281.7563, 281.8552, 281.9541, 282.0532, 282.1521, 282.251, 282.3499, 
    282.4487, 282.5479, 282.6467, 282.7456, 282.8445, 282.9421, 282.9529, 
    282.9639, 282.9746, 282.9854, 282.9961, 283.0068, 283.0176, 283.0283, 
    283.0391, 283.0498, 283.0605, 283.0713, 283.082, 283.019, 282.9214, 
    282.8237, 282.7261, 282.6284, 282.531, 282.4333, 282.3357, 282.238, 
    282.1404, 282.0427, 281.9451, 281.8474, 281.7654, 281.7124, 281.6594, 
    281.6067, 281.5537, 281.5007, 281.4478, 281.3948, 281.342, 281.2891, 
    281.2361, 281.1831, 281.1301, 281.0781, 281.0828, 281.0874, 281.092, 
    281.0969, 281.1016, 281.1062, 281.1108, 281.1155, 281.1201, 281.1248, 
    281.1294, 281.134, 281.1387, 281.1294, 281.1133, 281.0972, 281.0811, 
    281.0652, 281.0491, 281.033, 281.0171, 281.001, 280.9849, 280.9688, 
    280.9529, 280.9368, 280.9138, 280.8779, 280.842, 280.8062, 280.7705, 
    280.7346, 280.6987, 280.6628, 280.627, 280.5911, 280.5554, 280.5195, 
    280.4836, 280.4487, 280.468, 280.4875, 280.5068, 280.5261, 280.5457, 
    280.5649, 280.5845, 280.6038, 280.6233, 280.6426, 280.6619, 280.6814, 
    280.7007, 280.6978, 280.6843, 280.6711, 280.6577, 280.6443, 280.6309, 
    280.6177, 280.6042, 280.5908, 280.5774, 280.5642, 280.5508, 280.5374, 
    280.5149, 280.4753, 280.4355, 280.396, 280.3564, 280.3167, 280.2771, 
    280.2375, 280.1978, 280.1582, 280.1187, 280.0789, 280.0393, 279.9995, 
    279.9495, 279.8997, 279.8496, 279.7996, 279.7495, 279.6997, 279.6497, 
    279.5996, 279.5496, 279.4998, 279.4497, 279.3997, 279.3496, 279.283, 
    279.2087, 279.1343, 279.0598, 278.9856, 278.9111, 278.8367,
  278.0396, 278.0552, 278.071, 278.0867, 278.1025, 278.1182, 278.134, 
    278.1497, 278.1655, 278.1812, 278.197, 278.2126, 278.2527, 278.3386, 
    278.4248, 278.5107, 278.5967, 278.6829, 278.7688, 278.8547, 278.9409, 
    279.0269, 279.1128, 279.1987, 279.2849, 279.3721, 279.5591, 279.7461, 
    279.9331, 280.1201, 280.3071, 280.4941, 280.6812, 280.8682, 281.0552, 
    281.2422, 281.4292, 281.6162, 281.8032, 281.8457, 281.8198, 281.7937, 
    281.7676, 281.7417, 281.7156, 281.6897, 281.6636, 281.6377, 281.6116, 
    281.5857, 281.5596, 281.5334, 281.5442, 281.624, 281.7039, 281.7837, 
    281.8635, 281.9436, 282.0234, 282.1033, 282.1831, 282.2632, 282.343, 
    282.4229, 282.5027, 282.5852, 282.8665, 283.1479, 283.4292, 283.7107, 
    283.9919, 284.2732, 284.5547, 284.8359, 285.1174, 285.3987, 285.6802, 
    285.9614, 286.2429, 286.2012, 286.0066, 285.812, 285.6174, 285.4229, 
    285.2283, 285.0337, 284.8391, 284.6445, 284.45, 284.2554, 284.0608, 
    283.8662, 283.7415, 283.7488, 283.7561, 283.7634, 283.771, 283.7783, 
    283.7856, 283.793, 283.8003, 283.8079, 283.8152, 283.8225, 283.8298, 
    283.8372, 283.8323, 283.8271, 283.821, 283.8142, 283.8064, 283.7971, 
    283.7864, 283.7734, 283.7576, 283.738, 283.7129, 283.6799, 283.634, 
    283.2764, 282.905, 282.6318, 282.4224, 282.2568, 282.1223, 282.0112, 
    281.918, 281.8384, 281.7695, 281.7097, 281.657, 281.6104, 281.6194, 
    281.7251, 281.8308, 281.9363, 282.042, 282.1477, 282.2534, 282.3589, 
    282.4646, 282.5703, 282.676, 282.7817, 282.8872, 282.9915, 282.991, 
    282.9905, 282.9897, 282.9893, 282.9888, 282.9883, 282.9878, 282.9871, 
    282.9866, 282.9861, 282.9856, 282.9851, 282.9844, 282.9221, 282.8311, 
    282.7397, 282.6487, 282.5576, 282.4663, 282.3752, 282.2839, 282.1929, 
    282.1016, 282.0105, 281.9192, 281.8281, 281.7495, 281.6941, 281.6387, 
    281.5833, 281.5278, 281.4724, 281.417, 281.3616, 281.3064, 281.251, 
    281.1956, 281.1401, 281.0847, 281.0303, 281.0337, 281.0369, 281.0403, 
    281.0437, 281.0469, 281.0503, 281.0535, 281.0569, 281.0603, 281.0635, 
    281.0669, 281.0703, 281.0735, 281.0674, 281.0569, 281.0464, 281.0359, 
    281.0254, 281.0149, 281.0042, 280.9937, 280.9832, 280.9727, 280.9622, 
    280.9517, 280.9412, 280.9224, 280.8887, 280.8547, 280.821, 280.7874, 
    280.7534, 280.7197, 280.6858, 280.6521, 280.6182, 280.5845, 280.5508, 
    280.5168, 280.4839, 280.5032, 280.5225, 280.5417, 280.5613, 280.5806, 
    280.5999, 280.6191, 280.6384, 280.6577, 280.677, 280.6963, 280.7156, 
    280.7349, 280.7292, 280.7119, 280.6946, 280.677, 280.6597, 280.6423, 
    280.625, 280.6077, 280.5903, 280.573, 280.5557, 280.5381, 280.5208, 
    280.4978, 280.4639, 280.4302, 280.3962, 280.3625, 280.3286, 280.2949, 
    280.261, 280.2273, 280.1934, 280.1597, 280.1257, 280.092, 280.0579, 
    280.0076, 279.9573, 279.907, 279.8564, 279.8062, 279.7559, 279.7056, 
    279.655, 279.6047, 279.5544, 279.5042, 279.4539, 279.4033, 279.3337, 
    279.2554, 279.1768, 279.0984, 279.0198, 278.9414, 278.8628,
  278.281, 278.2981, 278.3152, 278.3323, 278.3494, 278.3665, 278.3835, 
    278.4006, 278.418, 278.4351, 278.4521, 278.4692, 278.5002, 278.5583, 
    278.6162, 278.6743, 278.7322, 278.7903, 278.8481, 278.9062, 278.9641, 
    279.0222, 279.0801, 279.1382, 279.196, 279.2556, 279.4485, 279.6411, 
    279.834, 280.0269, 280.2195, 280.4124, 280.6052, 280.7979, 280.9907, 
    281.1836, 281.3762, 281.5691, 281.762, 281.8167, 281.8059, 281.7952, 
    281.7842, 281.7734, 281.7627, 281.752, 281.7412, 281.7305, 281.7195, 
    281.7087, 281.698, 281.6873, 281.7097, 281.7954, 281.8809, 281.9666, 
    282.0522, 282.1377, 282.2234, 282.3088, 282.3945, 282.4802, 282.5657, 
    282.6514, 282.7371, 282.8245, 283.0605, 283.2966, 283.5327, 283.769, 
    284.0051, 284.2412, 284.4773, 284.7134, 284.9497, 285.1858, 285.4219, 
    285.658, 285.8943, 285.8579, 285.6929, 285.5276, 285.3625, 285.1975, 
    285.0325, 284.8672, 284.7021, 284.5371, 284.3718, 284.2068, 284.0417, 
    283.8767, 283.7759, 283.7966, 283.8176, 283.8384, 283.8594, 283.8801, 
    283.9011, 283.9219, 283.9429, 283.9636, 283.9846, 284.0054, 284.0264, 
    284.0469, 284.0386, 284.0295, 284.0193, 284.0081, 283.9956, 283.9812, 
    283.9651, 283.9465, 283.925, 283.8999, 283.8699, 283.8335, 283.7888, 
    283.5107, 283.1912, 282.9304, 282.7131, 282.5295, 282.3723, 282.2361, 
    282.1172, 282.0122, 281.9189, 281.8354, 281.7605, 281.6926, 281.688, 
    281.7925, 281.897, 282.0015, 282.106, 282.2104, 282.3149, 282.4194, 
    282.5239, 282.6284, 282.7332, 282.8376, 282.9421, 283.0449, 283.033, 
    283.021, 283.009, 282.9973, 282.9854, 282.9734, 282.9614, 282.9495, 
    282.9375, 282.9255, 282.9136, 282.9016, 282.8896, 282.8293, 282.7461, 
    282.6628, 282.5796, 282.4963, 282.4131, 282.3301, 282.2468, 282.1636, 
    282.0803, 281.9971, 281.9138, 281.8308, 281.7568, 281.7004, 281.644, 
    281.5876, 281.5312, 281.4749, 281.4185, 281.3621, 281.3057, 281.2493, 
    281.1929, 281.1365, 281.0801, 281.0247, 281.0237, 281.0229, 281.022, 
    281.0212, 281.0203, 281.0193, 281.0186, 281.0176, 281.0168, 281.0159, 
    281.0149, 281.0142, 281.0132, 281.01, 281.0056, 281.0012, 280.9968, 
    280.9924, 280.988, 280.9836, 280.979, 280.9746, 280.9702, 280.9658, 
    280.9614, 280.957, 280.9426, 280.9094, 280.8762, 280.843, 280.8098, 
    280.7764, 280.7432, 280.71, 280.6768, 280.6436, 280.6104, 280.5771, 
    280.5439, 280.5115, 280.5295, 280.5476, 280.5654, 280.5835, 280.6016, 
    280.6196, 280.6377, 280.6558, 280.6738, 280.6919, 280.7097, 280.7278, 
    280.7458, 280.7356, 280.7119, 280.6882, 280.6648, 280.6411, 280.6174, 
    280.594, 280.5703, 280.5466, 280.5232, 280.4995, 280.4761, 280.4524, 
    280.4285, 280.4036, 280.3789, 280.3542, 280.3296, 280.3047, 280.28, 
    280.2554, 280.2307, 280.2058, 280.1812, 280.1565, 280.1318, 280.1067, 
    280.0566, 280.0066, 279.9565, 279.9065, 279.8564, 279.8064, 279.7563, 
    279.7063, 279.6562, 279.6062, 279.5562, 279.5061, 279.4561, 279.3894, 
    279.3152, 279.241, 279.1665, 279.0923, 279.0178, 278.9436,
  278.5225, 278.541, 278.5593, 278.5779, 278.5964, 278.6147, 278.6333, 
    278.6519, 278.6702, 278.6887, 278.7073, 278.7256, 278.748, 278.7781, 
    278.8079, 278.8379, 278.8679, 278.8977, 278.9277, 278.9578, 278.9875, 
    279.0176, 279.0476, 279.0774, 279.1074, 279.1392, 279.3379, 279.5364, 
    279.7349, 279.9336, 280.1321, 280.3306, 280.5291, 280.7278, 280.9263, 
    281.1248, 281.3235, 281.522, 281.7205, 281.7876, 281.792, 281.7964, 
    281.8008, 281.8054, 281.8098, 281.8142, 281.8186, 281.8232, 281.8276, 
    281.832, 281.8364, 281.8408, 281.8752, 281.9668, 282.0581, 282.1494, 
    282.2407, 282.332, 282.4233, 282.5146, 282.606, 282.6973, 282.7886, 
    282.8799, 282.9712, 283.0637, 283.2546, 283.4456, 283.6365, 283.8274, 
    284.0183, 284.2092, 284.4001, 284.5911, 284.782, 284.9729, 285.1636, 
    285.3545, 285.5454, 285.5146, 285.3792, 285.2434, 285.1079, 284.9722, 
    284.8364, 284.7009, 284.5652, 284.4297, 284.2939, 284.1584, 284.0227, 
    283.887, 283.8103, 283.8447, 283.8789, 283.9133, 283.9478, 283.9822, 
    284.0166, 284.051, 284.0852, 284.1196, 284.1541, 284.1885, 284.2229, 
    284.2566, 284.2412, 284.2244, 284.2063, 284.1865, 284.1648, 284.1411, 
    284.1147, 284.0857, 284.0535, 284.0171, 283.9761, 283.9294, 283.8757, 
    283.6479, 283.3757, 283.1379, 282.9285, 282.7424, 282.5762, 282.4268, 
    282.2917, 282.1692, 282.0574, 281.9548, 281.8606, 281.7737, 281.7563, 
    281.8599, 281.9631, 282.0664, 282.1699, 282.2732, 282.3767, 282.48, 
    282.5833, 282.6868, 282.79, 282.8936, 282.9968, 283.0984, 283.0752, 
    283.0518, 283.0283, 283.0051, 282.9817, 282.9585, 282.9351, 282.9116, 
    282.8884, 282.865, 282.8416, 282.8184, 282.7949, 282.7363, 282.6611, 
    282.5857, 282.5105, 282.4353, 282.3601, 282.2849, 282.2095, 282.1343, 
    282.0591, 281.9839, 281.9084, 281.8333, 281.7642, 281.7068, 281.6494, 
    281.592, 281.5347, 281.4773, 281.4199, 281.3625, 281.3052, 281.2478, 
    281.1904, 281.1331, 281.0757, 281.019, 281.0139, 281.0088, 281.0037, 
    280.9988, 280.9937, 280.9885, 280.9834, 280.9783, 280.9731, 280.9683, 
    280.9631, 280.958, 280.9529, 280.9524, 280.9541, 280.9558, 280.9575, 
    280.9592, 280.9609, 280.9629, 280.9646, 280.9663, 280.968, 280.9697, 
    280.9714, 280.9731, 280.9629, 280.9302, 280.8975, 280.8647, 280.8323, 
    280.7996, 280.7668, 280.7341, 280.7014, 280.6687, 280.6362, 280.6035, 
    280.5708, 280.5388, 280.5557, 280.5725, 280.5891, 280.606, 280.6228, 
    280.6394, 280.6562, 280.6731, 280.6897, 280.7065, 280.7234, 280.74, 
    280.7568, 280.7417, 280.7119, 280.6821, 280.6523, 280.6226, 280.5928, 
    280.5627, 280.533, 280.5032, 280.4734, 280.4436, 280.4138, 280.3838, 
    280.3591, 280.3435, 280.3279, 280.312, 280.2964, 280.2808, 280.2651, 
    280.2495, 280.2339, 280.2183, 280.2026, 280.187, 280.1714, 280.1553, 
    280.1055, 280.0557, 280.0061, 279.9563, 279.9065, 279.8569, 279.8071, 
    279.7573, 279.7078, 279.658, 279.6082, 279.5586, 279.5088, 279.4451, 
    279.375, 279.3049, 279.2349, 279.1646, 279.0945, 279.0244,
  278.7642, 278.7839, 278.8037, 278.8235, 278.8433, 278.863, 278.8831, 
    278.9028, 278.9226, 278.9424, 278.9622, 278.9822, 278.9956, 278.9976, 
    278.9995, 279.0015, 279.0034, 279.0054, 279.0073, 279.009, 279.011, 
    279.0129, 279.0149, 279.0168, 279.0188, 279.0229, 279.2273, 279.4316, 
    279.636, 279.8401, 280.0444, 280.2488, 280.4531, 280.6575, 280.8618, 
    281.0662, 281.2705, 281.4749, 281.6792, 281.7583, 281.7781, 281.7979, 
    281.8174, 281.8372, 281.8567, 281.8765, 281.8962, 281.9158, 281.9355, 
    281.9553, 281.9749, 281.9946, 282.041, 282.1379, 282.2351, 282.332, 
    282.4292, 282.5261, 282.623, 282.7202, 282.8171, 282.9143, 283.0112, 
    283.1084, 283.2053, 283.303, 283.4485, 283.5942, 283.74, 283.8857, 
    284.0312, 284.177, 284.3228, 284.4685, 284.614, 284.7598, 284.9055, 
    285.0513, 285.1968, 285.1716, 285.0654, 284.9592, 284.853, 284.7468, 
    284.6406, 284.5344, 284.4285, 284.3223, 284.2161, 284.1099, 284.0037, 
    283.8975, 283.8447, 283.8926, 283.9404, 283.9883, 284.0361, 284.084, 
    284.1321, 284.1799, 284.2278, 284.2756, 284.3235, 284.3713, 284.4192, 
    284.4663, 284.4399, 284.4121, 284.3826, 284.3508, 284.3171, 284.2808, 
    284.2419, 284.2002, 284.155, 284.106, 284.053, 283.9951, 283.9316, 
    283.7383, 283.5046, 283.2908, 283.0942, 282.9133, 282.7458, 282.5906, 
    282.4463, 282.3118, 282.186, 282.0684, 281.958, 281.854, 281.825, 
    281.9272, 282.0293, 282.1316, 282.2339, 282.3359, 282.4382, 282.5405, 
    282.6428, 282.7449, 282.8472, 282.9495, 283.0515, 283.1519, 283.1172, 
    283.0825, 283.0476, 283.0129, 282.9783, 282.9434, 282.9087, 282.874, 
    282.8391, 282.8044, 282.7698, 282.7351, 282.7002, 282.6433, 282.5762, 
    282.5088, 282.4414, 282.3743, 282.3069, 282.2395, 282.1724, 282.105, 
    282.0378, 281.9705, 281.9031, 281.8359, 281.7717, 281.7134, 281.655, 
    281.5964, 281.5381, 281.4797, 281.4214, 281.363, 281.3047, 281.2461, 
    281.1877, 281.1294, 281.071, 281.0134, 281.0042, 280.9949, 280.9856, 
    280.9763, 280.9668, 280.9575, 280.9482, 280.939, 280.9297, 280.9204, 
    280.9111, 280.9019, 280.8926, 280.895, 280.9028, 280.9106, 280.9185, 
    280.9263, 280.9341, 280.9421, 280.95, 280.9578, 280.9656, 280.9734, 
    280.9812, 280.989, 280.9832, 280.9509, 280.9187, 280.8867, 280.8545, 
    280.8225, 280.7903, 280.7583, 280.7261, 280.6941, 280.6619, 280.6299, 
    280.5977, 280.5664, 280.582, 280.5974, 280.6128, 280.6284, 280.6438, 
    280.6594, 280.6748, 280.6904, 280.7058, 280.7214, 280.7368, 280.7524, 
    280.7678, 280.748, 280.7122, 280.676, 280.6399, 280.6038, 280.5679, 
    280.5317, 280.4956, 280.4597, 280.4236, 280.3875, 280.3516, 280.3154, 
    280.2898, 280.2832, 280.2766, 280.27, 280.2634, 280.2568, 280.2505, 
    280.2439, 280.2373, 280.2307, 280.2241, 280.2178, 280.2112, 280.2039, 
    280.1545, 280.105, 280.0557, 280.0061, 279.9568, 279.9075, 279.8579, 
    279.8086, 279.759, 279.7097, 279.6604, 279.6108, 279.5615, 279.5007, 
    279.4348, 279.3689, 279.303, 279.2371, 279.1711, 279.1052,
  279.0056, 279.0269, 279.0479, 279.0691, 279.0903, 279.1113, 279.1326, 
    279.1538, 279.175, 279.196, 279.2173, 279.2385, 279.2434, 279.2173, 
    279.1912, 279.165, 279.1389, 279.1128, 279.0867, 279.0605, 279.0344, 
    279.0083, 278.9822, 278.9561, 278.9299, 278.9065, 279.1167, 279.3267, 
    279.5369, 279.7468, 279.957, 280.1672, 280.3772, 280.5874, 280.7974, 
    281.0076, 281.2178, 281.4277, 281.6379, 281.7292, 281.7642, 281.7991, 
    281.834, 281.8689, 281.9038, 281.9387, 281.9736, 282.0085, 282.0435, 
    282.0784, 282.1135, 282.1484, 282.2065, 282.3093, 282.4121, 282.5149, 
    282.6177, 282.7202, 282.823, 282.9258, 283.0286, 283.1313, 283.2341, 
    283.3367, 283.4395, 283.5422, 283.6426, 283.7432, 283.8435, 283.9441, 
    284.0444, 284.145, 284.2454, 284.3459, 284.4463, 284.5469, 284.6472, 
    284.7478, 284.8481, 284.8284, 284.7517, 284.675, 284.5981, 284.5215, 
    284.4448, 284.3682, 284.2915, 284.2148, 284.1382, 284.0613, 283.9846, 
    283.908, 283.8792, 283.9404, 284.002, 284.0632, 284.1245, 284.186, 
    284.2473, 284.3088, 284.3701, 284.4316, 284.4929, 284.5544, 284.6157, 
    284.6758, 284.6355, 284.5933, 284.5491, 284.5029, 284.4548, 284.4043, 
    284.3513, 284.2957, 284.2373, 284.1758, 284.1111, 284.0427, 283.9705, 
    283.802, 283.5996, 283.4077, 283.2258, 283.0532, 282.8892, 282.7329, 
    282.584, 282.4419, 282.3062, 282.1765, 282.0522, 281.9333, 281.8936, 
    281.9946, 282.0957, 282.1968, 282.2979, 282.3989, 282.5, 282.6011, 
    282.7021, 282.8032, 282.9043, 283.0054, 283.1064, 283.2053, 283.1592, 
    283.113, 283.0669, 283.0208, 282.9746, 282.9285, 282.8823, 282.8362, 
    282.79, 282.7439, 282.6978, 282.6516, 282.6055, 282.5503, 282.491, 
    282.4316, 282.3723, 282.313, 282.2537, 282.1943, 282.135, 282.0757, 
    282.0164, 281.957, 281.8977, 281.8384, 281.7791, 281.7197, 281.6604, 
    281.6011, 281.5415, 281.4822, 281.4229, 281.3635, 281.304, 281.2446, 
    281.1853, 281.126, 281.0664, 281.0078, 280.9944, 280.9807, 280.9673, 
    280.9539, 280.9402, 280.9268, 280.9133, 280.8997, 280.8862, 280.8728, 
    280.8591, 280.8457, 280.8323, 280.8374, 280.8513, 280.8655, 280.8794, 
    280.8933, 280.9072, 280.9214, 280.9353, 280.9492, 280.9631, 280.9773, 
    280.9912, 281.0051, 281.0032, 280.9717, 280.9402, 280.9087, 280.877, 
    280.8455, 280.814, 280.7825, 280.751, 280.7192, 280.6877, 280.6562, 
    280.6248, 280.594, 280.6082, 280.6223, 280.6365, 280.6509, 280.665, 
    280.6792, 280.6934, 280.7078, 280.7219, 280.7361, 280.7502, 280.7646, 
    280.7788, 280.7544, 280.7122, 280.6699, 280.6274, 280.5852, 280.543, 
    280.5007, 280.4585, 280.416, 280.3738, 280.3315, 280.2893, 280.2468, 
    280.2202, 280.2229, 280.2253, 280.228, 280.2305, 280.2332, 280.2356, 
    280.238, 280.2407, 280.2432, 280.2458, 280.2483, 280.2507, 280.2524, 
    280.2034, 280.1543, 280.1052, 280.0562, 280.0071, 279.958, 279.9087, 
    279.8596, 279.8105, 279.7615, 279.7124, 279.6633, 279.6143, 279.5564, 
    279.4946, 279.4329, 279.3713, 279.3096, 279.2478, 279.186,
  279.2471, 279.2695, 279.2922, 279.3147, 279.3372, 279.3599, 279.3823, 
    279.4048, 279.4272, 279.45, 279.4724, 279.4949, 279.491, 279.437, 
    279.3828, 279.3286, 279.2744, 279.2205, 279.1663, 279.1121, 279.0579, 
    279.0037, 278.9497, 278.8955, 278.8413, 278.79, 279.0061, 279.2219, 
    279.4377, 279.6536, 279.8696, 280.0854, 280.3013, 280.5171, 280.7332, 
    280.949, 281.1648, 281.3806, 281.5967, 281.7002, 281.7502, 281.8003, 
    281.8506, 281.9006, 281.9509, 282.001, 282.0513, 282.1013, 282.1516, 
    282.2017, 282.252, 282.302, 282.3723, 282.4807, 282.5891, 282.6978, 
    282.8062, 282.9146, 283.0229, 283.1313, 283.24, 283.3484, 283.4568, 
    283.5652, 283.6736, 283.7815, 283.8367, 283.8918, 283.9473, 284.0024, 
    284.0576, 284.1128, 284.168, 284.2234, 284.2786, 284.3337, 284.3889, 
    284.4443, 284.4995, 284.4851, 284.438, 284.3906, 284.3435, 284.2961, 
    284.249, 284.2019, 284.1545, 284.1074, 284.0601, 284.0129, 283.9656, 
    283.9185, 283.9136, 283.9883, 284.0632, 284.1382, 284.2131, 284.2878, 
    284.3628, 284.4377, 284.5127, 284.5876, 284.6624, 284.7373, 284.8123, 
    284.8855, 284.8274, 284.7678, 284.7068, 284.644, 284.5798, 284.5139, 
    284.4463, 284.3767, 284.3054, 284.2319, 284.1565, 284.0789, 283.999, 
    283.8496, 283.6724, 283.5002, 283.333, 283.1702, 283.0117, 282.8574, 
    282.7073, 282.561, 282.4185, 282.2795, 282.144, 282.012, 281.9619, 
    282.0618, 282.1619, 282.2617, 282.3616, 282.4617, 282.5615, 282.6614, 
    282.7615, 282.8613, 282.9612, 283.0613, 283.1611, 283.2588, 283.2014, 
    283.1438, 283.0862, 283.0286, 282.9712, 282.9136, 282.856, 282.7986, 
    282.741, 282.6833, 282.626, 282.5684, 282.5107, 282.4575, 282.406, 
    282.3547, 282.3035, 282.252, 282.2007, 282.1492, 282.0979, 282.0466, 
    281.9951, 281.9438, 281.8923, 281.8411, 281.7866, 281.7261, 281.6658, 
    281.6055, 281.5449, 281.4846, 281.4243, 281.3638, 281.3035, 281.2432, 
    281.1826, 281.1223, 281.062, 281.0022, 280.9844, 280.9668, 280.949, 
    280.9314, 280.9136, 280.8958, 280.8782, 280.8604, 280.8428, 280.825, 
    280.8074, 280.7896, 280.7717, 280.7798, 280.8, 280.8201, 280.8403, 
    280.8604, 280.8804, 280.9006, 280.9207, 280.9407, 280.9609, 280.981, 
    281.001, 281.0212, 281.0234, 280.9924, 280.9614, 280.9304, 280.8994, 
    280.8687, 280.8376, 280.8066, 280.7756, 280.7446, 280.7136, 280.6826, 
    280.6516, 280.6213, 280.6343, 280.6472, 280.6602, 280.6731, 280.686, 
    280.699, 280.7122, 280.7251, 280.738, 280.751, 280.7639, 280.7769, 
    280.7898, 280.7607, 280.7122, 280.6636, 280.6152, 280.5667, 280.5181, 
    280.4695, 280.4211, 280.3726, 280.324, 280.2754, 280.2271, 280.1785, 
    280.1509, 280.1626, 280.1743, 280.1858, 280.1975, 280.2092, 280.2207, 
    280.2324, 280.2439, 280.2556, 280.2673, 280.2788, 280.2905, 280.301, 
    280.2524, 280.2036, 280.1548, 280.106, 280.0571, 280.0083, 279.9597, 
    279.9109, 279.8621, 279.8132, 279.7644, 279.7156, 279.667, 279.6121, 
    279.5544, 279.4971, 279.4395, 279.3818, 279.3245, 279.2668,
  279.4885, 279.5125, 279.5364, 279.5603, 279.5842, 279.6082, 279.6318, 
    279.6558, 279.6797, 279.7036, 279.7275, 279.7515, 279.7388, 279.6565, 
    279.5745, 279.4922, 279.4102, 279.3279, 279.2456, 279.1636, 279.0813, 
    278.999, 278.917, 278.8347, 278.7527, 278.6738, 278.8955, 279.1172, 
    279.3386, 279.5603, 279.782, 280.0037, 280.2253, 280.447, 280.6687, 
    280.8904, 281.1121, 281.3335, 281.5552, 281.6709, 281.7363, 281.8018, 
    281.8672, 281.9326, 281.998, 282.0632, 282.1287, 282.1941, 282.2595, 
    282.325, 282.3904, 282.4558, 282.5378, 282.6521, 282.7664, 282.8804, 
    282.9946, 283.1086, 283.2229, 283.3372, 283.4512, 283.5654, 283.6794, 
    283.7937, 283.9077, 284.0208, 284.0308, 284.0408, 284.0508, 284.0608, 
    284.0708, 284.0808, 284.0908, 284.1008, 284.1108, 284.1208, 284.1309, 
    284.1409, 284.1509, 284.1418, 284.1243, 284.1064, 284.0886, 284.071, 
    284.0532, 284.0354, 284.0176, 284, 283.9822, 283.9644, 283.9465, 283.929, 
    283.9478, 284.0364, 284.1248, 284.2131, 284.3015, 284.3899, 284.4783, 
    284.5667, 284.655, 284.7434, 284.832, 284.9204, 285.0088, 285.095, 
    285.0159, 284.9365, 284.8562, 284.7756, 284.6941, 284.6123, 284.5295, 
    284.4465, 284.3625, 284.2781, 284.1931, 284.1074, 284.021, 283.8862, 
    283.7302, 283.5754, 283.4219, 283.2693, 283.1179, 282.9678, 282.8186, 
    282.6707, 282.5237, 282.3779, 282.2332, 282.0894, 282.0305, 282.1292, 
    282.228, 282.3269, 282.4255, 282.5244, 282.6233, 282.7219, 282.8208, 
    282.9194, 283.0183, 283.1172, 283.2158, 283.3123, 283.2434, 283.1743, 
    283.1055, 283.0366, 282.9675, 282.8987, 282.8298, 282.7607, 282.6919, 
    282.6228, 282.554, 282.4851, 282.416, 282.3645, 282.321, 282.2776, 
    282.2344, 282.1909, 282.1475, 282.104, 282.0608, 282.0173, 281.9739, 
    281.9304, 281.887, 281.8438, 281.7939, 281.7327, 281.6711, 281.6099, 
    281.5483, 281.4871, 281.4258, 281.3643, 281.303, 281.2415, 281.1802, 
    281.1187, 281.0574, 280.9966, 280.9746, 280.9526, 280.9307, 280.9089, 
    280.887, 280.865, 280.843, 280.821, 280.7991, 280.7773, 280.7554, 
    280.7334, 280.7114, 280.7224, 280.7485, 280.7749, 280.801, 280.8274, 
    280.8535, 280.8799, 280.906, 280.9324, 280.9585, 280.9846, 281.011, 
    281.0371, 281.0437, 281.0132, 280.9829, 280.9524, 280.9219, 280.8916, 
    280.8611, 280.8308, 280.8003, 280.7698, 280.7395, 280.709, 280.6787, 
    280.6489, 280.6606, 280.6724, 280.6838, 280.6956, 280.7073, 280.719, 
    280.7307, 280.7424, 280.7539, 280.7656, 280.7773, 280.7891, 280.8008, 
    280.7671, 280.7122, 280.6575, 280.6028, 280.5481, 280.4932, 280.4385, 
    280.3838, 280.3291, 280.2742, 280.2195, 280.1648, 280.1099, 280.0815, 
    280.1023, 280.123, 280.1438, 280.1646, 280.1853, 280.2058, 280.2266, 
    280.2473, 280.2681, 280.2888, 280.3096, 280.3303, 280.3499, 280.3013, 
    280.2529, 280.2043, 280.1558, 280.1074, 280.0588, 280.0105, 279.9619, 
    279.9136, 279.865, 279.8167, 279.7681, 279.7195, 279.6677, 279.6145, 
    279.561, 279.5078, 279.4543, 279.4009, 279.3477,
  279.6484, 279.6792, 279.71, 279.7407, 279.7715, 279.802, 279.8328, 
    279.8635, 279.8943, 279.925, 279.9558, 279.9866, 279.978, 279.8943, 
    279.8108, 279.7271, 279.6436, 279.5598, 279.4763, 279.3926, 279.3091, 
    279.2253, 279.1418, 279.0581, 278.9746, 278.8943, 279.1038, 279.3132, 
    279.5229, 279.7324, 279.9421, 280.1516, 280.3611, 280.5708, 280.7803, 
    280.99, 281.1995, 281.4089, 281.6187, 281.7305, 281.7957, 281.8611, 
    281.9265, 281.9917, 282.0571, 282.1226, 282.1877, 282.2532, 282.3186, 
    282.384, 282.4492, 282.5146, 282.5903, 282.6858, 282.7815, 282.877, 
    282.9724, 283.0681, 283.1636, 283.259, 283.3547, 283.4502, 283.5457, 
    283.6414, 283.7368, 283.8311, 283.8281, 283.825, 283.8218, 283.8188, 
    283.8157, 283.8125, 283.8093, 283.8064, 283.8032, 283.8, 283.7971, 
    283.7939, 283.7908, 283.792, 283.7954, 283.7986, 283.8018, 283.8052, 
    283.8083, 283.8115, 283.8149, 283.8181, 283.8213, 283.8247, 283.8279, 
    283.8311, 283.8679, 283.9678, 284.0674, 284.1672, 284.2671, 284.3669, 
    284.4668, 284.5667, 284.6665, 284.7664, 284.8662, 284.9658, 285.0657, 
    285.1633, 285.083, 285.0022, 284.9204, 284.8379, 284.7546, 284.6704, 
    284.5852, 284.4995, 284.4126, 284.325, 284.2363, 284.1467, 284.0564, 
    283.9221, 283.769, 283.6174, 283.4673, 283.3188, 283.1719, 283.0264, 
    282.8823, 282.7397, 282.5984, 282.4587, 282.3203, 282.1831, 282.126, 
    282.2173, 282.3086, 282.3999, 282.4912, 282.5823, 282.6736, 282.7649, 
    282.8562, 282.9475, 283.0388, 283.1301, 283.2214, 283.3103, 283.238, 
    283.166, 283.0938, 283.0215, 282.9492, 282.877, 282.8049, 282.7327, 
    282.6604, 282.5881, 282.5161, 282.4438, 282.3716, 282.3218, 282.2825, 
    282.2434, 282.2041, 282.1648, 282.1255, 282.0864, 282.0471, 282.0078, 
    281.9685, 281.9292, 281.8901, 281.8508, 281.8044, 281.7451, 281.6855, 
    281.626, 281.5664, 281.5071, 281.4475, 281.3879, 281.3286, 281.269, 
    281.2095, 281.1501, 281.0906, 281.0315, 281.0061, 280.9805, 280.9548, 
    280.9294, 280.9038, 280.8782, 280.8528, 280.8271, 280.8015, 280.7761, 
    280.7505, 280.7249, 280.6995, 280.7107, 280.739, 280.7673, 280.7959, 
    280.8242, 280.8525, 280.8809, 280.9094, 280.9377, 280.9661, 280.9946, 
    281.0229, 281.0513, 281.0603, 281.0327, 281.0054, 280.9778, 280.9504, 
    280.9231, 280.8955, 280.8682, 280.8406, 280.8132, 280.7856, 280.7583, 
    280.731, 280.7041, 280.7131, 280.7222, 280.7312, 280.7402, 280.7493, 
    280.7583, 280.7673, 280.7764, 280.7854, 280.7944, 280.8035, 280.8125, 
    280.8215, 280.7864, 280.7305, 280.6746, 280.6187, 280.5627, 280.5068, 
    280.4512, 280.3953, 280.3394, 280.2834, 280.2275, 280.1716, 280.1157, 
    280.0864, 280.1064, 280.1265, 280.1465, 280.1665, 280.1865, 280.2065, 
    280.2263, 280.2463, 280.2664, 280.2864, 280.3064, 280.3264, 280.3452, 
    280.2961, 280.2473, 280.1985, 280.1494, 280.1006, 280.0515, 280.0027, 
    279.9536, 279.9048, 279.8557, 279.8069, 279.7581, 279.709, 279.6599, 
    279.6111, 279.562, 279.5129, 279.4639, 279.415, 279.366,
  279.7468, 279.7886, 279.8303, 279.8721, 279.9138, 279.9556, 279.9973, 
    280.0388, 280.0806, 280.1223, 280.1641, 280.2058, 280.2107, 280.1458, 
    280.0806, 280.0154, 279.9504, 279.8853, 279.8201, 279.7551, 279.6899, 
    279.6248, 279.5598, 279.4946, 279.4294, 279.3672, 279.5513, 279.7354, 
    279.9194, 280.1035, 280.2876, 280.4717, 280.6558, 280.8401, 281.0242, 
    281.2083, 281.3923, 281.5764, 281.7605, 281.8562, 281.9102, 281.9639, 
    282.0178, 282.0715, 282.1255, 282.1794, 282.2332, 282.2871, 282.3408, 
    282.3948, 282.4485, 282.5024, 282.5579, 282.6167, 282.6753, 282.7339, 
    282.7925, 282.8513, 282.9099, 282.9685, 283.0273, 283.0859, 283.1445, 
    283.2031, 283.262, 283.3201, 283.3279, 283.3357, 283.3435, 283.3516, 
    283.3594, 283.3672, 283.3752, 283.3831, 283.3909, 283.3989, 283.4067, 
    283.4146, 283.4224, 283.4373, 283.4551, 283.4731, 283.491, 283.5088, 
    283.5269, 283.5447, 283.5627, 283.5806, 283.5986, 283.6165, 283.6345, 
    283.6523, 283.7019, 283.8118, 283.9214, 284.031, 284.1409, 284.2505, 
    284.3601, 284.4697, 284.5796, 284.6892, 284.7988, 284.9084, 285.0183, 
    285.1257, 285.0605, 284.9937, 284.925, 284.8542, 285.0134, 284.9973, 
    284.9827, 284.9695, 284.9573, 284.946, 284.9355, 284.926, 284.917, 
    283.9697, 283.8054, 283.646, 283.4917, 283.342, 283.1968, 283.0559, 
    282.9189, 282.7861, 282.6567, 282.5312, 282.4092, 282.2903, 282.2417, 
    282.3208, 282.3999, 282.4788, 282.5579, 282.6367, 282.7158, 282.7949, 
    282.8738, 282.9529, 283.0317, 283.1108, 283.1897, 283.2668, 283.1973, 
    283.1279, 283.0586, 282.9893, 282.9199, 282.8506, 282.781, 282.7117, 
    282.6423, 282.573, 282.5037, 282.4343, 282.3647, 282.3169, 282.2788, 
    282.241, 282.2029, 282.165, 282.127, 282.0891, 282.0513, 282.0132, 
    281.9753, 281.9373, 281.8994, 281.8613, 281.8174, 281.762, 281.7065, 
    281.6511, 281.5957, 281.54, 281.4846, 281.4292, 281.3738, 281.3184, 
    281.2629, 281.2075, 281.1521, 281.0972, 281.0684, 281.0396, 281.011, 
    280.9822, 280.9534, 280.9246, 280.896, 280.8672, 280.8384, 280.8096, 
    280.781, 280.7522, 280.7234, 280.7332, 280.7607, 280.7883, 280.8159, 
    280.8435, 280.8711, 280.8987, 280.9263, 280.9539, 280.9814, 281.009, 
    281.0366, 281.0642, 281.0742, 281.0515, 281.0288, 281.0061, 280.9834, 
    280.9607, 280.938, 280.9153, 280.8928, 280.8701, 280.8474, 280.8247, 
    280.802, 280.7798, 280.7852, 280.7905, 280.7959, 280.8015, 280.8069, 
    280.8123, 280.8176, 280.823, 280.8284, 280.8337, 280.8391, 280.8447, 
    280.8501, 280.8154, 280.7622, 280.709, 280.656, 280.6028, 280.5496, 
    280.4963, 280.4434, 280.3901, 280.3369, 280.2837, 280.2307, 280.1775, 
    280.147, 280.1589, 280.1709, 280.1829, 280.1946, 280.2065, 280.2185, 
    280.2305, 280.2422, 280.2542, 280.2661, 280.2781, 280.2898, 280.3008, 
    280.2507, 280.2007, 280.1509, 280.1008, 280.0508, 280.0007, 279.9509, 
    279.9009, 279.8508, 279.801, 279.751, 279.7009, 279.6509, 279.6047, 
    279.5601, 279.5156, 279.4709, 279.4265, 279.3818, 279.3374,
  279.8452, 279.8979, 279.9507, 280.0034, 280.0562, 280.1089, 280.1616, 
    280.2144, 280.2671, 280.3196, 280.3723, 280.425, 280.4436, 280.397, 
    280.3503, 280.304, 280.2573, 280.2107, 280.1641, 280.1174, 280.0708, 
    280.0242, 279.9775, 279.9312, 279.8845, 279.8401, 279.9988, 280.1575, 
    280.3159, 280.4746, 280.6333, 280.792, 280.9504, 281.1091, 281.2678, 
    281.4265, 281.585, 281.7437, 281.9023, 281.9822, 282.0244, 282.0669, 
    282.1091, 282.1516, 282.1938, 282.2361, 282.2786, 282.3208, 282.3633, 
    282.4055, 282.448, 282.4902, 282.5254, 282.5474, 282.5691, 282.5908, 
    282.6125, 282.6345, 282.6562, 282.678, 282.7, 282.7217, 282.7434, 
    282.7651, 282.7871, 282.8088, 282.8276, 282.8464, 282.8655, 282.8843, 
    282.9031, 282.9219, 282.9409, 282.9597, 282.9785, 282.9976, 283.0164, 
    283.0352, 283.054, 283.0823, 283.115, 283.1475, 283.1802, 283.2126, 
    283.2454, 283.2778, 283.3105, 283.343, 283.3757, 283.4082, 283.4409, 
    283.4736, 283.5361, 283.6558, 283.7754, 283.8948, 284.0144, 284.134, 
    284.2534, 284.373, 284.4924, 284.6121, 284.7317, 284.8511, 284.9707, 
    285.0881, 285.0376, 284.9851, 284.9299, 284.8721, 285.1255, 285.1301, 
    285.134, 285.1375, 285.1404, 285.1431, 285.1455, 285.1479, 285.1499, 
    284.0315, 283.8513, 283.6814, 283.521, 283.3694, 283.2256, 283.0891, 
    282.9597, 282.8364, 282.7192, 282.6074, 282.5005, 282.3987, 282.3577, 
    282.4243, 282.491, 282.5579, 282.6245, 282.6912, 282.7581, 282.8247, 
    282.8914, 282.958, 283.0249, 283.0916, 283.1582, 283.2231, 283.1565, 
    283.0901, 283.0234, 282.957, 282.8904, 282.824, 282.7573, 282.6909, 
    282.6243, 282.5579, 282.4912, 282.4246, 282.3582, 282.312, 282.2751, 
    282.2385, 282.2019, 282.1653, 282.1287, 282.0918, 282.0552, 282.0186, 
    281.9819, 281.9453, 281.9084, 281.8718, 281.8301, 281.7788, 281.7273, 
    281.676, 281.6248, 281.5732, 281.522, 281.4705, 281.4192, 281.3679, 
    281.3164, 281.2651, 281.2136, 281.1626, 281.1306, 281.0989, 281.0669, 
    281.0349, 281.0029, 280.9709, 280.9392, 280.9072, 280.8752, 280.8433, 
    280.8113, 280.7795, 280.7476, 280.7556, 280.7825, 280.8091, 280.8359, 
    280.8628, 280.8894, 280.9163, 280.9431, 280.9697, 280.9966, 281.0234, 
    281.05, 281.0769, 281.0881, 281.0701, 281.0522, 281.0344, 281.0164, 
    280.9985, 280.9807, 280.9626, 280.9448, 280.927, 280.9089, 280.8911, 
    280.8733, 280.8557, 280.8574, 280.8591, 280.8608, 280.8625, 280.8643, 
    280.8662, 280.8679, 280.8696, 280.8713, 280.873, 280.875, 280.8767, 
    280.8784, 280.8445, 280.7939, 280.7437, 280.6931, 280.6426, 280.5923, 
    280.5417, 280.4912, 280.4409, 280.3904, 280.3398, 280.2896, 280.239, 
    280.2075, 280.2114, 280.2151, 280.219, 280.2229, 280.2266, 280.2305, 
    280.2344, 280.238, 280.2419, 280.2456, 280.2495, 280.2534, 280.2563, 
    280.2053, 280.1543, 280.1033, 280.0522, 280.0012, 279.9502, 279.8992, 
    279.8481, 279.7971, 279.7461, 279.6951, 279.644, 279.593, 279.5493, 
    279.5093, 279.4692, 279.4292, 279.3889, 279.3489, 279.3088,
  279.9438, 280.0076, 280.071, 280.1348, 280.1985, 280.2622, 280.3259, 
    280.3896, 280.4534, 280.5171, 280.5806, 280.6443, 280.6765, 280.6484, 
    280.6204, 280.5923, 280.5642, 280.5361, 280.5081, 280.4797, 280.4517, 
    280.4236, 280.3955, 280.3674, 280.3394, 280.313, 280.4463, 280.5793, 
    280.7126, 280.8457, 280.979, 281.1121, 281.2451, 281.3784, 281.5115, 
    281.6448, 281.7778, 281.9111, 282.0442, 282.1079, 282.1389, 282.1697, 
    282.2004, 282.2314, 282.2622, 282.293, 282.3237, 282.3547, 282.3855, 
    282.4163, 282.4473, 282.478, 282.4929, 282.478, 282.4629, 282.4478, 
    282.4326, 282.4177, 282.4026, 282.3875, 282.3723, 282.3574, 282.3423, 
    282.3271, 282.312, 282.2976, 282.3274, 282.3572, 282.3872, 282.417, 
    282.4468, 282.4768, 282.5066, 282.5364, 282.5662, 282.5962, 282.626, 
    282.6558, 282.6858, 282.7273, 282.7747, 282.822, 282.8691, 282.9165, 
    282.9639, 283.011, 283.0583, 283.1055, 283.1528, 283.2002, 283.2473, 
    283.2947, 283.3704, 283.4998, 283.6292, 283.7585, 283.8879, 284.0173, 
    284.1467, 284.2761, 284.4055, 284.5349, 284.6643, 284.7937, 284.9231, 
    285.0505, 285.0144, 284.9758, 284.9348, 284.8911, 285.2107, 285.2273, 
    285.2415, 285.2537, 285.2642, 285.2737, 285.282, 285.2893, 285.2959, 
    284.1152, 283.9116, 283.7263, 283.5571, 283.4021, 283.2593, 283.1272, 
    283.0051, 282.8916, 282.7859, 282.6873, 282.5947, 282.5083, 282.4734, 
    282.5278, 282.5823, 282.6367, 282.6912, 282.7456, 282.8, 282.8545, 
    282.9089, 282.9634, 283.0178, 283.0723, 283.1267, 283.1794, 283.116, 
    283.0522, 282.9885, 282.9248, 282.8611, 282.7974, 282.7336, 282.6699, 
    282.6062, 282.5425, 282.4788, 282.415, 282.3513, 282.3069, 282.2715, 
    282.2363, 282.2009, 282.1655, 282.1301, 282.0947, 282.0593, 282.0239, 
    281.9885, 281.9531, 281.9177, 281.8826, 281.843, 281.7957, 281.7483, 
    281.7009, 281.6538, 281.6064, 281.5591, 281.5117, 281.4646, 281.4172, 
    281.3699, 281.3225, 281.2754, 281.2283, 281.1931, 281.158, 281.1228, 
    281.0876, 281.0525, 281.0173, 280.9824, 280.9473, 280.9121, 280.877, 
    280.8418, 280.8066, 280.7717, 280.7781, 280.8042, 280.8301, 280.856, 
    280.8821, 280.908, 280.9338, 280.9597, 280.9858, 281.0117, 281.0376, 
    281.0637, 281.0896, 281.1018, 281.0889, 281.0757, 281.0625, 281.0493, 
    281.0364, 281.0232, 281.01, 280.9968, 280.9836, 280.9707, 280.9575, 
    280.9443, 280.9314, 280.9294, 280.9277, 280.9258, 280.9238, 280.9219, 
    280.9202, 280.9182, 280.9163, 280.9143, 280.9124, 280.9106, 280.9087, 
    280.9067, 280.8735, 280.8259, 280.7781, 280.7302, 280.6826, 280.6348, 
    280.5872, 280.5393, 280.4917, 280.4438, 280.396, 280.3484, 280.3005, 
    280.2681, 280.2639, 280.2595, 280.2554, 280.251, 280.2468, 280.2424, 
    280.2383, 280.2339, 280.2297, 280.2253, 280.2212, 280.2168, 280.2117, 
    280.1597, 280.1077, 280.0557, 280.0034, 279.9514, 279.8994, 279.8474, 
    279.7952, 279.7432, 279.6912, 279.6392, 279.5869, 279.5349, 279.4941, 
    279.4585, 279.4229, 279.3872, 279.3516, 279.3159, 279.2803,
  280.0422, 280.1169, 280.1917, 280.2664, 280.3408, 280.4155, 280.4902, 
    280.5649, 280.6396, 280.7144, 280.7891, 280.8635, 280.9094, 280.8997, 
    280.8901, 280.8806, 280.8711, 280.8613, 280.8518, 280.8423, 280.8328, 
    280.823, 280.8135, 280.804, 280.7944, 280.7861, 280.8938, 281.0015, 
    281.1091, 281.2168, 281.3245, 281.4321, 281.5398, 281.6477, 281.7554, 
    281.863, 281.9707, 282.0784, 282.186, 282.2339, 282.2532, 282.2725, 
    282.2917, 282.3113, 282.3306, 282.3499, 282.3691, 282.3884, 282.408, 
    282.4272, 282.4465, 282.4658, 282.4607, 282.4087, 282.3567, 282.3047, 
    282.2527, 282.2009, 282.1489, 282.0969, 282.0449, 281.9932, 281.9412, 
    281.8892, 281.8372, 281.7864, 281.8271, 281.8682, 281.9089, 281.9497, 
    281.9905, 282.0315, 282.0723, 282.113, 282.1541, 282.1948, 282.2356, 
    282.2764, 282.3174, 282.3726, 282.4343, 282.4963, 282.5583, 282.6204, 
    282.6821, 282.7441, 282.8062, 282.8682, 282.9299, 282.9919, 283.054, 
    283.116, 283.2046, 283.3438, 283.4832, 283.6223, 283.7615, 283.9009, 
    284.04, 284.1794, 284.3186, 284.458, 284.5972, 284.7363, 284.8757, 
    285.0129, 284.9907, 284.9666, 284.9402, 284.9116, 285.2771, 285.3015, 
    285.3215, 285.3389, 285.3535, 285.3662, 285.3774, 285.3875, 285.3962, 
    284.2344, 283.9939, 283.7854, 283.603, 283.4421, 283.2991, 283.1711, 
    283.0562, 282.9521, 282.8574, 282.771, 282.6919, 282.6189, 282.5891, 
    282.6313, 282.6736, 282.7156, 282.7578, 282.8, 282.8423, 282.8843, 
    282.9265, 282.9688, 283.011, 283.053, 283.0952, 283.136, 283.0752, 
    283.0142, 282.9534, 282.8926, 282.8315, 282.7708, 282.71, 282.6489, 
    282.5881, 282.5273, 282.4663, 282.4055, 282.3447, 282.302, 282.2678, 
    282.2339, 282.1997, 282.1658, 282.1316, 282.0974, 282.0635, 282.0293, 
    281.9954, 281.9612, 281.927, 281.8931, 281.8557, 281.8125, 281.7693, 
    281.7261, 281.6829, 281.6396, 281.5962, 281.553, 281.5098, 281.4666, 
    281.4233, 281.3801, 281.3369, 281.2937, 281.2554, 281.217, 281.1787, 
    281.1404, 281.1021, 281.064, 281.0256, 280.9873, 280.949, 280.9106, 
    280.8723, 280.834, 280.7957, 280.8005, 280.8257, 280.8508, 280.876, 
    280.9011, 280.9263, 280.9514, 280.9766, 281.0017, 281.0269, 281.052, 
    281.0771, 281.1023, 281.1157, 281.1074, 281.0991, 281.0908, 281.0823, 
    281.074, 281.0657, 281.0574, 281.0491, 281.0405, 281.0322, 281.0239, 
    281.0156, 281.0073, 281.0017, 280.9961, 280.9905, 280.9851, 280.9795, 
    280.9739, 280.9685, 280.9629, 280.9573, 280.9519, 280.9463, 280.9407, 
    280.9353, 280.9026, 280.8577, 280.8125, 280.7676, 280.7224, 280.6775, 
    280.6323, 280.5874, 280.5425, 280.4973, 280.4524, 280.4072, 280.3623, 
    280.3286, 280.3162, 280.304, 280.2915, 280.2793, 280.2668, 280.2544, 
    280.2422, 280.2297, 280.2173, 280.2051, 280.1926, 280.1804, 280.1672, 
    280.1143, 280.061, 280.0081, 279.9548, 279.9019, 279.8486, 279.7957, 
    279.7424, 279.6892, 279.6362, 279.583, 279.53, 279.4768, 279.4387, 
    279.4077, 279.3765, 279.3452, 279.3142, 279.283, 279.2517,
  280.1406, 280.2263, 280.312, 280.3977, 280.4834, 280.5688, 280.6545, 
    280.7402, 280.8259, 280.9116, 280.9973, 281.083, 281.1421, 281.1511, 
    281.1599, 281.1689, 281.178, 281.1868, 281.1958, 281.2046, 281.2136, 
    281.2224, 281.2314, 281.2402, 281.2493, 281.259, 281.3413, 281.4233, 
    281.5056, 281.5879, 281.6702, 281.7524, 281.8345, 281.9167, 281.999, 
    282.0813, 282.1636, 282.2456, 282.3279, 282.3596, 282.3674, 282.3755, 
    282.3833, 282.3911, 282.3989, 282.4067, 282.4146, 282.4224, 282.4302, 
    282.438, 282.4458, 282.4536, 282.4282, 282.3394, 282.2505, 282.1616, 
    282.0728, 281.9841, 281.8953, 281.8064, 281.7175, 281.6289, 281.54, 
    281.4512, 281.3623, 281.2751, 281.3271, 281.3789, 281.4307, 281.4824, 
    281.5344, 281.5862, 281.6379, 281.6897, 281.7417, 281.7935, 281.8452, 
    281.897, 281.949, 282.0176, 282.0942, 282.1709, 282.2473, 282.324, 
    282.4006, 282.4773, 282.554, 282.6306, 282.7073, 282.7837, 282.8604, 
    282.937, 283.0388, 283.1877, 283.3369, 283.4861, 283.6353, 283.7844, 
    283.9333, 284.0825, 284.2317, 284.3809, 284.53, 284.679, 284.8281, 
    284.9751, 284.9666, 284.9568, 284.946, 284.9341, 285.3308, 285.3599, 
    285.3838, 285.4041, 285.4209, 285.4355, 285.4482, 285.4595, 285.4692, 
    284.4182, 284.1128, 283.866, 283.6626, 283.4922, 283.3474, 283.2224, 
    283.114, 283.0188, 282.9343, 282.8594, 282.792, 282.7312, 282.7048, 
    282.7349, 282.7646, 282.7947, 282.8245, 282.8545, 282.8843, 282.9143, 
    282.9441, 282.9741, 283.0039, 283.0339, 283.0637, 283.0923, 283.0344, 
    282.9763, 282.9182, 282.8604, 282.8022, 282.7441, 282.686, 282.6282, 
    282.5701, 282.512, 282.4539, 282.396, 282.3379, 282.2971, 282.2642, 
    282.2314, 282.1987, 282.1658, 282.1331, 282.1003, 282.0676, 282.0347, 
    282.002, 281.9692, 281.9363, 281.9036, 281.8687, 281.8293, 281.7903, 
    281.751, 281.7119, 281.6726, 281.6335, 281.5942, 281.5552, 281.5159, 
    281.4768, 281.4377, 281.3984, 281.3591, 281.3176, 281.2761, 281.2349, 
    281.1934, 281.1519, 281.1104, 281.0688, 281.0273, 280.9858, 280.9443, 
    280.9028, 280.8613, 280.8198, 280.8232, 280.8474, 280.8718, 280.8962, 
    280.9204, 280.9448, 280.9692, 280.9934, 281.0178, 281.0422, 281.0664, 
    281.0908, 281.1152, 281.1296, 281.1262, 281.1226, 281.1189, 281.1155, 
    281.1118, 281.1082, 281.1045, 281.1011, 281.0974, 281.0938, 281.0903, 
    281.0867, 281.083, 281.0737, 281.0647, 281.0554, 281.0461, 281.0371, 
    281.0278, 281.0188, 281.0095, 281.0002, 280.9912, 280.9819, 280.9727, 
    280.9636, 280.9316, 280.8894, 280.8472, 280.8047, 280.7625, 280.7202, 
    280.6777, 280.6355, 280.593, 280.5508, 280.5085, 280.4661, 280.4238, 
    280.3892, 280.3687, 280.3481, 280.3279, 280.3074, 280.2869, 280.2664, 
    280.2461, 280.2256, 280.2051, 280.1848, 280.1643, 280.1438, 280.1228, 
    280.0686, 280.0144, 279.9604, 279.9062, 279.8521, 279.7979, 279.7437, 
    279.6897, 279.6355, 279.5813, 279.5271, 279.4731, 279.4189, 279.3835, 
    279.3567, 279.3301, 279.3035, 279.2766, 279.25, 279.2231,
  280.239, 280.3357, 280.4324, 280.5291, 280.6257, 280.7224, 280.8191, 
    280.9155, 281.0122, 281.1089, 281.2056, 281.3022, 281.375, 281.4023, 
    281.4299, 281.4573, 281.4849, 281.5122, 281.5396, 281.5671, 281.5945, 
    281.6218, 281.6494, 281.6768, 281.7041, 281.7319, 281.7888, 281.8455, 
    281.9023, 281.959, 282.0156, 282.0725, 282.1292, 282.186, 282.2427, 
    282.2996, 282.3562, 282.4131, 282.4697, 282.4856, 282.4819, 282.4783, 
    282.4746, 282.4709, 282.4673, 282.4636, 282.46, 282.4561, 282.4524, 
    282.4487, 282.4451, 282.4414, 282.3958, 282.27, 282.1443, 282.0186, 
    281.8931, 281.7673, 281.6416, 281.5159, 281.3901, 281.2646, 281.1389, 
    281.0132, 280.8875, 280.7642, 280.8269, 280.8896, 280.9524, 281.0154, 
    281.0781, 281.1409, 281.2036, 281.2666, 281.3293, 281.3921, 281.4548, 
    281.5178, 281.5806, 281.6626, 281.7539, 281.8452, 281.9365, 282.0278, 
    282.1191, 282.2104, 282.3018, 282.3931, 282.4844, 282.5757, 282.667, 
    282.7583, 282.8728, 283.032, 283.1909, 283.3499, 283.5088, 283.6677, 
    283.8267, 283.9858, 284.1448, 284.3037, 284.4626, 284.6216, 284.7805, 
    284.9375, 284.9419, 284.9465, 284.9521, 284.9583, 285.3748, 285.4072, 
    285.4336, 285.4553, 285.4736, 285.4893, 285.5027, 285.5146, 285.5249, 
    284.7393, 284.2998, 283.9832, 283.7439, 283.5569, 283.4065, 283.2832, 
    283.1799, 283.0925, 283.0173, 282.9521, 282.895, 282.8445, 282.8208, 
    282.8384, 282.856, 282.8735, 282.8911, 282.9089, 282.9265, 282.9441, 
    282.9617, 282.9792, 282.9971, 283.0146, 283.0322, 283.0488, 282.9937, 
    282.9385, 282.8833, 282.8279, 282.7727, 282.7175, 282.6624, 282.6072, 
    282.552, 282.4968, 282.4417, 282.3865, 282.3311, 282.292, 282.2605, 
    282.229, 282.1975, 282.166, 282.1345, 282.103, 282.0715, 282.04, 
    282.0085, 281.9771, 281.9456, 281.9141, 281.8813, 281.8462, 281.811, 
    281.7761, 281.741, 281.7058, 281.6707, 281.6355, 281.6006, 281.5654, 
    281.5303, 281.4951, 281.46, 281.4248, 281.3801, 281.3354, 281.2908, 
    281.2461, 281.2014, 281.1567, 281.1121, 281.0674, 281.0227, 280.978, 
    280.9331, 280.8884, 280.8438, 280.8457, 280.8691, 280.8928, 280.9163, 
    280.9397, 280.9634, 280.9868, 281.0103, 281.0337, 281.0574, 281.0808, 
    281.1042, 281.1279, 281.1436, 281.1448, 281.146, 281.1472, 281.1484, 
    281.1497, 281.1506, 281.1519, 281.1531, 281.1543, 281.1555, 281.1567, 
    281.158, 281.1589, 281.146, 281.1331, 281.1204, 281.1074, 281.0947, 
    281.0818, 281.0691, 281.0562, 281.0432, 281.0305, 281.0176, 281.0049, 
    280.9919, 280.9609, 280.9211, 280.8816, 280.842, 280.8022, 280.7627, 
    280.7231, 280.6836, 280.6438, 280.6042, 280.5647, 280.5251, 280.4854, 
    280.4497, 280.4211, 280.3926, 280.364, 280.3354, 280.3071, 280.2786, 
    280.25, 280.2214, 280.1929, 280.1643, 280.1357, 280.1072, 280.0784, 
    280.0232, 279.968, 279.9128, 279.8577, 279.8022, 279.7471, 279.6919, 
    279.6367, 279.5815, 279.5264, 279.4712, 279.416, 279.3608, 279.3281, 
    279.3059, 279.2837, 279.2615, 279.2393, 279.217, 279.1946,
  280.2483, 280.3567, 280.4651, 280.5737, 280.6821, 280.7905, 280.8989, 
    281.0073, 281.1157, 281.2241, 281.3325, 281.4409, 281.5273, 281.572, 
    281.6165, 281.6611, 281.7056, 281.75, 281.7947, 281.8391, 281.8838, 
    281.9282, 281.9727, 282.0173, 282.0618, 282.1064, 282.1465, 282.1868, 
    282.2268, 282.2671, 282.3071, 282.3474, 282.3877, 282.4277, 282.468, 
    282.5081, 282.5483, 282.5886, 282.6287, 282.6409, 282.6394, 282.6382, 
    282.637, 282.6355, 282.6343, 282.6331, 282.6316, 282.6304, 282.6292, 
    282.6279, 282.6265, 282.6252, 282.5737, 282.4272, 282.2805, 282.1338, 
    281.9871, 281.8406, 281.6938, 281.5471, 281.4006, 281.2539, 281.1072, 
    280.9607, 280.814, 280.6697, 280.7268, 280.7839, 280.8408, 280.8979, 
    280.9551, 281.012, 281.0691, 281.1262, 281.1831, 281.2402, 281.2974, 
    281.3542, 281.4114, 281.4954, 281.5923, 281.6892, 281.7859, 281.8828, 
    281.9797, 282.0767, 282.1733, 282.2703, 282.3672, 282.4639, 282.5608, 
    282.6577, 282.7756, 282.9338, 283.092, 283.2502, 283.4087, 283.5669, 
    283.7251, 283.8833, 284.0415, 284.1997, 284.3579, 284.5161, 284.6743, 
    284.8306, 284.8428, 284.8564, 284.8723, 284.8906, 285.4006, 285.4412, 
    285.4739, 285.501, 285.5234, 285.5427, 285.5591, 285.5735, 285.5862, 
    285.0354, 284.4932, 284.1311, 283.8726, 283.6785, 283.5273, 283.4065, 
    283.3074, 283.2251, 283.1553, 283.0955, 283.0435, 282.9983, 282.9727, 
    282.9761, 282.9795, 282.9829, 282.9863, 282.9897, 282.9932, 282.9968, 
    283.0002, 283.0037, 283.0071, 283.0105, 283.0139, 283.0166, 282.9692, 
    282.9216, 282.8743, 282.8267, 282.7793, 282.7317, 282.6843, 282.637, 
    282.5894, 282.542, 282.4944, 282.447, 282.3994, 282.3599, 282.3237, 
    282.2876, 282.2515, 282.2151, 282.179, 282.1428, 282.1067, 282.0706, 
    282.0344, 281.9983, 281.9622, 281.926, 281.8916, 281.8606, 281.8296, 
    281.7983, 281.7673, 281.7363, 281.7051, 281.6741, 281.6428, 281.6118, 
    281.5808, 281.5496, 281.5186, 281.4873, 281.4473, 281.407, 281.3669, 
    281.3269, 281.2869, 281.2466, 281.2065, 281.1665, 281.1265, 281.0862, 
    281.0461, 281.0061, 280.9661, 280.9688, 280.9915, 281.0139, 281.0366, 
    281.0593, 281.082, 281.1047, 281.1274, 281.1501, 281.1729, 281.1956, 
    281.2183, 281.2407, 281.2539, 281.249, 281.2441, 281.2395, 281.2346, 
    281.2297, 281.2249, 281.22, 281.2153, 281.2104, 281.2056, 281.2007, 
    281.1958, 281.1909, 281.1768, 281.1624, 281.1482, 281.134, 281.1196, 
    281.1055, 281.0913, 281.0771, 281.0627, 281.0486, 281.0344, 281.02, 
    281.0059, 280.9785, 280.9446, 280.9106, 280.876, 280.8413, 280.8062, 
    280.7708, 280.7349, 280.6987, 280.6624, 280.6255, 280.5884, 280.5508, 
    280.5151, 280.4836, 280.4519, 280.4204, 280.3889, 280.3574, 280.3259, 
    280.2944, 280.2629, 280.2312, 280.1997, 280.1682, 280.1367, 280.1047, 
    280.0493, 279.9937, 279.9382, 279.8828, 279.8271, 279.7717, 279.7163, 
    279.6606, 279.6052, 279.5496, 279.4941, 279.4387, 279.3831, 279.3489, 
    279.3247, 279.3008, 279.2769, 279.2534, 279.2302, 279.207,
  280.1826, 280.3035, 280.4243, 280.5452, 280.666, 280.7869, 280.9077, 
    281.0286, 281.1494, 281.2703, 281.3911, 281.512, 281.6121, 281.6726, 
    281.7329, 281.7935, 281.854, 281.9143, 281.9749, 282.0354, 282.0957, 
    282.1562, 282.2168, 282.2771, 282.3376, 282.3977, 282.4287, 282.46, 
    282.491, 282.5222, 282.5532, 282.5842, 282.6155, 282.6465, 282.6775, 
    282.7087, 282.7397, 282.771, 282.802, 282.8206, 282.8335, 282.8462, 
    282.8589, 282.8718, 282.8845, 282.8972, 282.9102, 282.9229, 282.9355, 
    282.9485, 282.9612, 282.9739, 282.9292, 282.7749, 282.6206, 282.4663, 
    282.312, 282.158, 282.0037, 281.8494, 281.6951, 281.541, 281.3867, 
    281.2324, 281.0781, 280.9263, 280.9634, 281.0007, 281.0378, 281.0752, 
    281.1123, 281.1494, 281.1868, 281.2239, 281.2612, 281.2983, 281.3354, 
    281.3728, 281.4099, 281.4863, 281.5811, 281.6758, 281.7705, 281.8652, 
    281.96, 282.0544, 282.1492, 282.2439, 282.3386, 282.4333, 282.5281, 
    282.6228, 282.7363, 282.8848, 283.0332, 283.1819, 283.3303, 283.4788, 
    283.6274, 283.7759, 283.9243, 284.073, 284.2214, 284.3701, 284.5186, 
    284.6653, 284.6814, 284.6995, 284.7202, 284.7444, 285.4158, 285.4692, 
    285.5122, 285.5479, 285.5774, 285.6028, 285.6245, 285.6436, 285.6602, 
    285.1343, 284.6155, 284.269, 284.0215, 283.8357, 283.6912, 283.5754, 
    283.481, 283.4019, 283.3352, 283.2778, 283.2283, 283.1848, 283.155, 
    283.1426, 283.1304, 283.1179, 283.1055, 283.0933, 283.0808, 283.0686, 
    283.0562, 283.0437, 283.0315, 283.019, 283.0066, 282.9939, 282.9583, 
    282.9229, 282.8872, 282.8516, 282.8159, 282.7803, 282.7446, 282.709, 
    282.6736, 282.6379, 282.6023, 282.5667, 282.531, 282.4885, 282.4429, 
    282.397, 282.3513, 282.3054, 282.2598, 282.2139, 282.1682, 282.1223, 
    282.0767, 282.0308, 281.9851, 281.9395, 281.9001, 281.8728, 281.8457, 
    281.8186, 281.7915, 281.7644, 281.7373, 281.71, 281.6829, 281.6558, 
    281.6287, 281.6016, 281.5742, 281.5471, 281.5183, 281.4893, 281.4602, 
    281.4314, 281.4023, 281.3733, 281.3445, 281.3154, 281.2864, 281.2576, 
    281.2285, 281.1995, 281.1707, 281.1763, 281.198, 281.22, 281.2417, 
    281.2634, 281.2854, 281.3071, 281.3291, 281.3508, 281.3726, 281.3945, 
    281.4163, 281.4382, 281.4453, 281.4255, 281.4055, 281.3855, 281.3657, 
    281.3457, 281.3257, 281.3057, 281.2859, 281.2659, 281.2458, 281.2261, 
    281.2061, 281.1863, 281.1724, 281.1587, 281.145, 281.1313, 281.1174, 
    281.1038, 281.0901, 281.0764, 281.0625, 281.0488, 281.0352, 281.0215, 
    281.0076, 280.9866, 280.9614, 280.9358, 280.9092, 280.8818, 280.854, 
    280.8252, 280.7954, 280.7649, 280.7334, 280.7009, 280.6675, 280.6331, 
    280.5994, 280.5693, 280.5396, 280.5095, 280.4795, 280.4495, 280.4194, 
    280.3896, 280.3596, 280.3296, 280.2996, 280.2695, 280.2397, 280.2092, 
    280.1541, 280.0989, 280.0437, 279.9885, 279.9333, 279.8782, 279.8232, 
    279.7681, 279.7129, 279.6577, 279.6025, 279.5474, 279.4922, 279.4504, 
    279.416, 279.3826, 279.3501, 279.3186, 279.2881, 279.2585,
  280.1167, 280.25, 280.3833, 280.5166, 280.6499, 280.7832, 280.9165, 
    281.0498, 281.1831, 281.3164, 281.4497, 281.583, 281.6968, 281.7732, 
    281.8496, 281.926, 282.0022, 282.0786, 282.155, 282.2314, 282.3079, 
    282.3843, 282.4607, 282.5369, 282.6133, 282.6892, 282.7112, 282.7332, 
    282.7551, 282.7771, 282.7991, 282.8213, 282.8433, 282.8652, 282.8872, 
    282.9092, 282.9312, 282.9534, 282.9753, 283.0005, 283.0273, 283.0542, 
    283.0811, 283.1079, 283.1348, 283.1616, 283.1885, 283.2153, 283.2422, 
    283.269, 283.2959, 283.3225, 283.2844, 283.1226, 282.9607, 282.7988, 
    282.637, 282.4753, 282.3135, 282.1516, 281.9897, 281.8279, 281.666, 
    281.5044, 281.3425, 281.1829, 281.2002, 281.2175, 281.2349, 281.2522, 
    281.2695, 281.2871, 281.3044, 281.3218, 281.3391, 281.3564, 281.3738, 
    281.3911, 281.4084, 281.4771, 281.5696, 281.6621, 281.7549, 281.8474, 
    281.9399, 282.0325, 282.1252, 282.2178, 282.3103, 282.4031, 282.4956, 
    282.5881, 282.6968, 282.8357, 282.9744, 283.1133, 283.2522, 283.3909, 
    283.5298, 283.6687, 283.8074, 283.9463, 284.0852, 284.2239, 284.3628, 
    284.5, 284.5198, 284.5425, 284.5681, 284.5981, 285.4309, 285.4971, 
    285.5505, 285.5945, 285.6316, 285.6628, 285.6899, 285.7134, 285.7339, 
    285.2332, 284.7375, 284.407, 284.1707, 283.9932, 283.855, 283.7446, 
    283.6543, 283.5789, 283.5151, 283.4604, 283.4131, 283.3716, 283.3374, 
    283.3093, 283.281, 283.2529, 283.2249, 283.1965, 283.1685, 283.1404, 
    283.1121, 283.084, 283.0557, 283.0276, 282.9995, 282.9714, 282.9475, 
    282.9238, 282.9001, 282.8765, 282.8525, 282.8289, 282.8052, 282.7812, 
    282.7576, 282.7339, 282.7102, 282.6863, 282.6626, 282.6172, 282.562, 
    282.5066, 282.4512, 282.3958, 282.3403, 282.2849, 282.2295, 282.1741, 
    282.1187, 282.0632, 282.0081, 281.9526, 281.9084, 281.8853, 281.8621, 
    281.8389, 281.8157, 281.7925, 281.7693, 281.7461, 281.7229, 281.6997, 
    281.6765, 281.6533, 281.6301, 281.6072, 281.5894, 281.5713, 281.5535, 
    281.5356, 281.5178, 281.5, 281.4822, 281.4644, 281.4465, 281.4287, 
    281.4109, 281.3931, 281.3752, 281.3838, 281.4048, 281.4258, 281.4468, 
    281.4678, 281.4885, 281.5095, 281.5305, 281.5515, 281.5725, 281.5935, 
    281.6145, 281.6355, 281.637, 281.6018, 281.5667, 281.5317, 281.4966, 
    281.4617, 281.4265, 281.3914, 281.3564, 281.3213, 281.2864, 281.2512, 
    281.2161, 281.1814, 281.1682, 281.155, 281.1418, 281.1287, 281.1152, 
    281.1021, 281.0889, 281.0757, 281.0625, 281.0491, 281.0359, 281.0227, 
    281.0095, 280.9949, 280.9788, 280.9622, 280.9446, 280.9263, 280.907, 
    280.8867, 280.8655, 280.843, 280.8193, 280.7942, 280.7678, 280.7397, 
    280.7107, 280.6829, 280.6548, 280.627, 280.5991, 280.571, 280.5432, 
    280.5151, 280.4873, 280.4595, 280.4314, 280.4036, 280.3755, 280.3472, 
    280.2925, 280.2378, 280.1831, 280.1284, 280.0737, 280.019, 279.9644, 
    279.9097, 279.855, 279.8003, 279.7456, 279.6909, 279.6362, 279.5825, 
    279.5317, 279.4839, 279.4385, 279.3958, 279.3552, 279.3167,
  280.0508, 280.1965, 280.3423, 280.488, 280.6338, 280.7795, 280.9253, 
    281.071, 281.2168, 281.3625, 281.5083, 281.6541, 281.7815, 281.8738, 
    281.9661, 282.0583, 282.1506, 282.2429, 282.3352, 282.4275, 282.5198, 
    282.6123, 282.7046, 282.7969, 282.8892, 282.9805, 282.9934, 283.0063, 
    283.0193, 283.0322, 283.0452, 283.0581, 283.071, 283.084, 283.0969, 
    283.1099, 283.1228, 283.1355, 283.1484, 283.1804, 283.2214, 283.2622, 
    283.3032, 283.344, 283.385, 283.4258, 283.4668, 283.5078, 283.5486, 
    283.5896, 283.6304, 283.6714, 283.6396, 283.4702, 283.3008, 283.1313, 
    282.9619, 282.7927, 282.6233, 282.4539, 282.2844, 282.115, 281.9456, 
    281.7761, 281.6067, 281.4392, 281.4368, 281.4343, 281.4319, 281.4294, 
    281.427, 281.4246, 281.4221, 281.4194, 281.417, 281.4146, 281.4121, 
    281.4097, 281.4072, 281.4678, 281.5583, 281.6487, 281.7393, 281.8296, 
    281.9202, 282.0105, 282.1011, 282.1917, 282.282, 282.3726, 282.4629, 
    282.5535, 282.6572, 282.7864, 282.9155, 283.0447, 283.1738, 283.303, 
    283.4321, 283.5613, 283.6904, 283.8196, 283.9487, 284.0779, 284.207, 
    284.3347, 284.3584, 284.3853, 284.416, 284.4519, 285.446, 285.5251, 
    285.5889, 285.6414, 285.6855, 285.7229, 285.7551, 285.7832, 285.8079, 
    285.7908, 285.751, 285.7058, 285.6536, 285.5925, 285.5203, 285.4336, 
    285.3279, 283.7559, 283.6951, 283.6428, 283.5979, 283.5583, 283.5198, 
    283.4758, 283.4319, 283.3879, 283.344, 283.3, 283.2561, 283.2122, 
    283.168, 283.124, 283.0801, 283.0361, 282.9922, 282.9487, 282.9368, 
    282.925, 282.9131, 282.9011, 282.8892, 282.8774, 282.8655, 282.8535, 
    282.8418, 282.8298, 282.8179, 282.8062, 282.7942, 282.7461, 282.6812, 
    282.616, 282.551, 282.4861, 282.4209, 282.356, 282.291, 282.2258, 
    282.1609, 282.0959, 282.0308, 281.9658, 281.9167, 281.8975, 281.8782, 
    281.8591, 281.8398, 281.8206, 281.8013, 281.7822, 281.7629, 281.7437, 
    281.7244, 281.7053, 281.686, 281.667, 281.6604, 281.6536, 281.647, 
    281.6401, 281.6335, 281.6267, 281.6201, 281.6133, 281.6067, 281.5999, 
    281.5933, 281.5864, 281.5798, 281.5913, 281.6113, 281.6316, 281.6516, 
    281.6719, 281.6919, 281.7119, 281.7322, 281.7522, 281.7725, 281.7925, 
    281.8125, 281.8328, 281.8284, 281.7781, 281.728, 281.6777, 281.6277, 
    281.5774, 281.5273, 281.4771, 281.427, 281.3767, 281.3267, 281.2764, 
    281.2263, 281.1768, 281.1641, 281.1514, 281.1387, 281.1257, 281.113, 
    281.1003, 281.0876, 281.075, 281.0623, 281.0496, 281.0366, 281.0239, 
    281.0112, 281.0029, 280.9966, 280.9897, 280.9824, 280.9746, 281.9644, 
    282.0481, 282.1201, 282.1829, 282.2378, 282.2864, 282.3296, 282.3684, 
    282.3926, 282.3958, 282.3987, 282.4016, 282.4048, 282.4077, 282.4106, 
    282.4138, 282.4167, 282.4199, 282.4229, 282.4258, 282.429, 282.4312, 
    282.3833, 282.3357, 282.2878, 282.2402, 282.1926, 282.1448, 282.0972, 
    282.0493, 282.0017, 281.9541, 281.9062, 281.8586, 281.8108, 281.7488, 
    281.6736, 281.5898, 281.4956, 281.3892, 281.2678, 279.3831,
  279.9851, 280.1433, 280.3015, 280.4595, 280.6177, 280.7759, 280.9341, 
    281.0923, 281.2505, 281.4087, 281.5669, 281.7251, 281.8662, 281.9744, 
    282.0825, 282.1909, 282.2991, 282.4072, 282.5154, 282.6238, 282.7319, 
    282.8401, 282.9485, 283.0566, 283.1648, 283.272, 283.2759, 283.2795, 
    283.2834, 283.2874, 283.291, 283.2949, 283.2988, 283.3027, 283.3064, 
    283.3103, 283.3142, 283.3179, 283.3218, 283.3604, 283.4153, 283.4702, 
    283.5251, 283.5803, 283.6353, 283.6902, 283.7451, 283.8, 283.8552, 
    283.9102, 283.9651, 284.02, 283.9949, 283.8179, 283.6409, 283.4639, 
    283.2869, 283.1101, 282.9331, 282.7561, 282.5791, 282.4021, 282.2251, 
    282.0481, 281.8711, 281.6958, 281.6736, 281.6511, 281.6289, 281.6067, 
    281.5842, 281.562, 281.5396, 281.5173, 281.4951, 281.4727, 281.4504, 
    281.428, 281.4058, 281.4585, 281.5469, 281.6353, 281.7236, 281.812, 
    281.9004, 281.9885, 282.0769, 282.1653, 282.2537, 282.342, 282.4304, 
    282.5188, 282.6177, 282.7373, 282.8567, 282.9761, 283.0957, 283.2151, 
    283.3345, 283.4539, 283.5735, 283.6929, 283.8123, 283.9316, 284.0513, 
    284.1694, 284.197, 284.2283, 284.2642, 284.3057, 285.4612, 285.553, 
    285.6272, 285.6882, 285.7395, 285.783, 285.8206, 285.853, 285.8816, 
    285.8669, 285.8293, 285.7861, 285.7366, 285.6785, 285.6099, 285.5276, 
    285.427, 283.9326, 283.875, 283.8254, 283.7825, 283.7449, 283.7021, 
    283.6423, 283.5825, 283.5229, 283.4631, 283.4033, 283.3435, 283.2839, 
    283.2241, 283.1643, 283.1045, 283.0447, 282.9851, 282.926, 282.926, 
    282.926, 282.926, 282.926, 282.926, 282.926, 282.9258, 282.9258, 
    282.9258, 282.9258, 282.9258, 282.9258, 282.9258, 282.8748, 282.8003, 
    282.7256, 282.6509, 282.5762, 282.5015, 282.427, 282.3523, 282.2776, 
    282.2029, 282.1284, 282.0537, 281.979, 281.925, 281.9097, 281.8945, 
    281.8792, 281.864, 281.8486, 281.8335, 281.8181, 281.803, 281.7876, 
    281.7725, 281.7571, 281.7419, 281.7268, 281.7312, 281.7358, 281.7402, 
    281.7446, 281.749, 281.7534, 281.7578, 281.7622, 281.7666, 281.771, 
    281.7754, 281.78, 281.7844, 281.7988, 281.8181, 281.8374, 281.8567, 
    281.876, 281.8953, 281.9146, 281.9338, 281.9529, 281.9722, 281.9915, 
    282.0107, 282.03, 282.0198, 281.9546, 281.8892, 281.824, 281.7588, 
    281.6934, 281.6282, 281.5627, 281.4976, 281.4324, 281.3669, 281.3018, 
    281.2366, 281.1721, 281.1599, 281.1475, 281.1353, 281.123, 281.1108, 
    281.0986, 281.0864, 281.0742, 281.062, 281.0498, 281.0376, 281.0254, 
    281.0129, 281.0115, 281.0149, 281.0188, 281.0229, 281.0276, 282.123, 
    282.2085, 282.2805, 282.3423, 282.3955, 282.4421, 282.4834, 282.5198, 
    282.5435, 282.5491, 282.5549, 282.5608, 282.5667, 282.5723, 282.5781, 
    282.584, 282.5898, 282.5955, 282.6013, 282.6072, 282.613, 282.6179, 
    282.5708, 282.5237, 282.4766, 282.4294, 282.3826, 282.3354, 282.2883, 
    282.2412, 282.1941, 282.147, 282.0999, 282.053, 282.0059, 281.9487, 
    281.8806, 281.8042, 281.7173, 281.6177, 281.5027, 279.4597,
  279.9192, 280.0898, 280.2605, 280.4312, 280.6018, 280.7725, 280.9429, 
    281.1135, 281.2842, 281.4548, 281.6255, 281.7961, 281.9507, 282.075, 
    282.199, 282.3232, 282.4475, 282.5715, 282.6958, 282.8198, 282.9441, 
    283.0681, 283.1924, 283.3164, 283.4407, 283.5632, 283.5581, 283.5527, 
    283.5476, 283.5422, 283.5371, 283.5317, 283.5266, 283.5212, 283.5161, 
    283.5107, 283.5056, 283.5002, 283.4951, 283.5403, 283.6091, 283.6782, 
    283.7473, 283.8164, 283.8855, 283.9543, 284.0234, 284.0925, 284.1616, 
    284.2307, 284.2998, 284.3687, 284.3503, 284.1658, 283.9812, 283.7966, 
    283.6121, 283.4272, 283.2427, 283.0581, 282.8735, 282.689, 282.5044, 
    282.3198, 282.1353, 281.9524, 281.9102, 281.8682, 281.8259, 281.7837, 
    281.7417, 281.6995, 281.6572, 281.6152, 281.573, 281.5308, 281.4888, 
    281.4465, 281.4043, 281.4495, 281.5356, 281.6218, 281.708, 281.7942, 
    281.8804, 281.9666, 282.053, 282.1392, 282.2253, 282.3115, 282.3977, 
    282.4839, 282.5784, 282.688, 282.7979, 282.9075, 283.0173, 283.1272, 
    283.2368, 283.3467, 283.4563, 283.5662, 283.676, 283.7856, 283.8955, 
    284.0042, 284.0354, 284.071, 284.1121, 284.1592, 285.4763, 285.5811, 
    285.6655, 285.7351, 285.7935, 285.843, 285.8857, 285.9229, 285.9556, 
    285.9431, 285.9075, 285.8667, 285.8196, 285.7644, 285.6995, 285.6216, 
    285.5261, 284.1096, 284.0549, 284.0081, 283.9673, 283.9316, 283.8845, 
    283.8088, 283.7334, 283.658, 283.5823, 283.5068, 283.4312, 283.3557, 
    283.28, 283.2046, 283.1289, 283.0535, 282.9778, 282.9036, 282.9153, 
    282.9272, 282.939, 282.9507, 282.9626, 282.9744, 282.9863, 282.998, 
    283.01, 283.0217, 283.0337, 283.0454, 283.0571, 283.0037, 282.9194, 
    282.835, 282.7507, 282.6665, 282.5823, 282.498, 282.4136, 282.3293, 
    282.2451, 282.1609, 282.0764, 281.9922, 281.9333, 281.9221, 281.9106, 
    281.8994, 281.8882, 281.877, 281.8655, 281.8542, 281.843, 281.8315, 
    281.8203, 281.8091, 281.7976, 281.7869, 281.8022, 281.8179, 281.8335, 
    281.8491, 281.8645, 281.8801, 281.8958, 281.9111, 281.9268, 281.9424, 
    281.9578, 281.9734, 281.989, 282.0063, 282.0249, 282.0432, 282.0618, 
    282.0801, 282.0984, 282.1169, 282.1353, 282.1538, 282.1721, 282.1904, 
    282.209, 282.2273, 282.2112, 282.1309, 282.0505, 281.9702, 281.8896, 
    281.8093, 281.729, 281.6484, 281.5681, 281.4878, 281.4075, 281.3269, 
    281.2466, 281.1672, 281.1555, 281.1438, 281.1321, 281.1204, 281.1086, 
    281.0969, 281.0852, 281.0735, 281.0618, 281.05, 281.0383, 281.0266, 
    281.0149, 281.02, 281.0339, 281.0496, 281.0667, 281.0862, 282.249, 
    282.3335, 282.4036, 282.4629, 282.5137, 282.5579, 282.5962, 282.6301, 
    282.6528, 282.6606, 282.6685, 282.6763, 282.6841, 282.6919, 282.6997, 
    282.7075, 282.7153, 282.7231, 282.731, 282.7388, 282.7466, 282.7534, 
    282.7068, 282.6602, 282.6135, 282.5669, 282.5203, 282.4736, 282.427, 
    282.3804, 282.3337, 282.2871, 282.2407, 282.1941, 282.1475, 282.0945, 
    282.033, 281.9631, 281.8831, 281.7908, 281.6829, 279.5491,
  279.8533, 280.0364, 280.2195, 280.4026, 280.5857, 280.7688, 280.9519, 
    281.1348, 281.3179, 281.501, 281.6841, 281.8672, 282.0354, 282.1755, 
    282.3157, 282.4558, 282.5957, 282.7358, 282.876, 283.0161, 283.156, 
    283.2961, 283.4363, 283.5764, 283.7163, 283.8547, 283.8403, 283.8262, 
    283.8118, 283.7974, 283.783, 283.7688, 283.7544, 283.74, 283.7256, 
    283.7114, 283.697, 283.6826, 283.6685, 283.72, 283.8032, 283.8862, 
    283.9695, 284.0525, 284.1357, 284.2188, 284.3018, 284.385, 284.468, 
    284.5513, 284.6343, 284.7175, 284.7056, 284.5134, 284.3213, 284.1292, 
    283.937, 283.7446, 283.5525, 283.3604, 283.1682, 282.9761, 282.7839, 
    282.5918, 282.3994, 282.209, 282.147, 282.085, 282.0229, 281.9609, 
    281.8989, 281.8369, 281.7749, 281.7129, 281.6509, 281.5889, 281.5269, 
    281.4648, 281.4028, 281.4402, 281.5242, 281.6084, 281.6924, 281.7764, 
    281.8606, 281.9446, 282.0288, 282.1128, 282.197, 282.281, 282.3652, 
    282.4492, 282.5388, 282.6389, 282.739, 282.8391, 282.9392, 283.0391, 
    283.1392, 283.2393, 283.3394, 283.4395, 283.5396, 283.6396, 283.7397, 
    283.8389, 283.874, 283.9141, 283.96, 284.0129, 285.4915, 285.6089, 
    285.7039, 285.782, 285.8474, 285.9031, 285.9512, 285.9927, 286.0293, 
    286.0195, 285.9856, 285.947, 285.9026, 285.8506, 285.7891, 285.7153, 
    285.6252, 284.2866, 284.2349, 284.1904, 284.1521, 284.1184, 284.0669, 
    283.9756, 283.8843, 283.7927, 283.7014, 283.6101, 283.5188, 283.4275, 
    283.3359, 283.2446, 283.1533, 283.062, 282.9707, 282.8809, 282.9045, 
    282.9282, 282.9519, 282.9756, 282.9993, 283.0229, 283.0466, 283.0703, 
    283.094, 283.1177, 283.1414, 283.165, 283.1887, 283.1323, 283.0386, 
    282.9446, 282.8506, 282.7568, 282.6628, 282.5688, 282.4751, 282.3811, 
    282.2871, 282.1934, 282.0994, 282.0054, 281.9417, 281.9343, 281.927, 
    281.9197, 281.9124, 281.905, 281.8977, 281.8904, 281.8828, 281.8755, 
    281.8682, 281.8608, 281.8535, 281.8467, 281.8733, 281.9001, 281.9268, 
    281.9534, 281.9802, 282.0068, 282.0334, 282.0601, 282.0869, 282.1135, 
    282.1401, 282.1667, 282.1936, 282.2141, 282.2314, 282.249, 282.2666, 
    282.2842, 282.3018, 282.3193, 282.3369, 282.3545, 282.3721, 282.3896, 
    282.407, 282.4246, 282.4028, 282.3071, 282.2117, 282.1162, 282.0208, 
    281.9253, 281.8298, 281.7341, 281.6387, 281.5432, 281.4478, 281.3523, 
    281.2568, 281.1626, 281.1514, 281.1401, 281.1289, 281.1177, 281.1064, 
    281.0952, 281.084, 281.0728, 281.0615, 281.0503, 281.0391, 281.0278, 
    281.0166, 281.0286, 281.0535, 281.0818, 281.114, 281.1511, 282.3513, 
    282.4333, 282.501, 282.5576, 282.6055, 282.647, 282.6826, 282.7141, 
    282.7358, 282.7454, 282.7546, 282.7639, 282.7732, 282.7827, 282.792, 
    282.8013, 282.8108, 282.8201, 282.8293, 282.8386, 282.8481, 282.8564, 
    282.8101, 282.7639, 282.7175, 282.6714, 282.625, 282.5789, 282.5325, 
    282.4861, 282.4399, 282.3936, 282.3474, 282.301, 282.2549, 282.2056, 
    282.1497, 282.0857, 282.0122, 281.9265, 281.8257, 279.6545,
  279.8721, 280.0605, 280.2488, 280.4373, 280.6255, 280.814, 281.0022, 
    281.1907, 281.3789, 281.5674, 281.7556, 281.9441, 282.1177, 282.2627, 
    282.408, 282.553, 282.6982, 282.8435, 282.9885, 283.1338, 283.2788, 
    283.4241, 283.5693, 283.7144, 283.8596, 284.0029, 283.9827, 283.9622, 
    283.9419, 283.9214, 283.9011, 283.8806, 283.8604, 283.8401, 283.8196, 
    283.7993, 283.7788, 283.7585, 283.738, 283.7891, 283.874, 283.9587, 
    284.0437, 284.1284, 284.2134, 284.2981, 284.3831, 284.4678, 284.5527, 
    284.6375, 284.7224, 284.8071, 284.802, 284.6257, 284.4495, 284.2732, 
    284.0972, 283.9209, 283.7446, 283.5684, 283.3923, 283.2161, 283.0398, 
    282.8635, 282.6875, 282.5125, 282.4343, 282.3562, 282.2781, 282.2002, 
    282.1221, 282.0439, 281.9658, 281.8879, 281.8098, 281.7317, 281.6536, 
    281.5757, 281.4976, 281.5234, 281.5989, 281.6741, 281.7493, 281.8245, 
    281.8997, 281.9751, 282.0503, 282.1255, 282.2007, 282.2759, 282.3513, 
    282.4265, 282.5078, 282.6011, 282.6951, 282.79, 282.8857, 282.9824, 
    283.0798, 283.1782, 283.2776, 283.3779, 283.479, 283.5811, 283.6841, 
    283.7871, 283.8274, 283.873, 283.925, 283.9854, 285.5925, 285.7068, 
    285.8018, 285.8816, 285.9497, 286.0085, 286.0598, 286.105, 286.145, 
    286.1365, 286.1035, 286.0659, 286.0234, 285.9744, 285.9172, 285.8501, 
    285.7698, 284.4146, 284.3601, 284.3132, 284.2727, 284.2371, 284.1794, 
    284.0742, 283.9702, 283.8672, 283.7651, 283.6638, 283.5635, 283.4641, 
    283.3655, 283.2681, 283.1711, 283.0752, 282.9802, 282.8877, 282.9119, 
    282.936, 282.9602, 282.9844, 283.0083, 283.0325, 283.0566, 283.0808, 
    283.105, 283.1292, 283.1533, 283.1775, 283.2017, 283.1445, 283.0493, 
    282.9541, 282.8591, 282.7639, 282.6687, 282.5737, 282.4785, 282.3833, 
    282.2881, 282.1931, 282.0979, 282.0027, 281.9392, 281.9353, 281.9312, 
    281.9272, 281.9231, 281.9189, 281.915, 281.9109, 281.907, 281.9028, 
    281.8987, 281.8948, 281.8906, 281.8872, 281.9199, 281.9529, 281.9858, 
    282.0186, 282.0515, 282.0845, 282.1174, 282.1501, 282.1831, 282.2161, 
    282.2488, 282.2817, 282.3147, 282.3347, 282.3489, 282.363, 282.3774, 
    282.3916, 282.4058, 282.4199, 282.4341, 282.4482, 282.4624, 282.4766, 
    282.491, 282.5051, 282.4797, 282.3811, 282.2825, 282.1836, 282.085, 
    281.9861, 281.8875, 281.7888, 281.6899, 281.5913, 281.4927, 281.3938, 
    281.2952, 281.1978, 281.1873, 281.1768, 281.1665, 281.156, 281.1455, 
    281.135, 281.1245, 281.114, 281.1035, 281.0933, 281.0828, 281.0723, 
    281.0618, 281.0769, 281.1069, 281.1414, 281.1809, 281.2271, 282.4187, 
    282.4983, 282.5637, 282.6179, 282.6638, 282.7034, 282.7375, 282.7676, 
    282.7888, 282.7998, 282.8108, 282.8218, 282.8328, 282.8438, 282.8547, 
    282.8657, 282.8767, 282.8877, 282.8987, 282.9097, 282.9207, 282.9307, 
    282.8853, 282.8398, 282.7947, 282.7493, 282.7039, 282.6587, 282.6133, 
    282.5679, 282.5227, 282.4773, 282.4319, 282.3867, 282.3413, 282.2935, 
    282.239, 282.177, 282.1052, 282.0212, 281.9224, 279.7183,
  279.9707, 280.1577, 280.3445, 280.5315, 280.7183, 280.9053, 281.092, 
    281.2791, 281.4658, 281.6526, 281.8396, 282.0264, 282.1973, 282.3372, 
    282.4773, 282.6174, 282.7573, 282.8975, 283.0374, 283.1775, 283.3176, 
    283.4575, 283.5977, 283.7375, 283.8777, 284.0159, 283.9924, 283.969, 
    283.9453, 283.9219, 283.8984, 283.8748, 283.8513, 283.8279, 283.8042, 
    283.7808, 283.7573, 283.7336, 283.7102, 283.7534, 283.8284, 283.9033, 
    283.9783, 284.0532, 284.1279, 284.2029, 284.2778, 284.3528, 284.4277, 
    284.5027, 284.5776, 284.6526, 284.6538, 284.5159, 284.3779, 284.2397, 
    284.1018, 283.9639, 283.8257, 283.6877, 283.5498, 283.4116, 283.2737, 
    283.1357, 282.9976, 282.8601, 282.7695, 282.679, 282.5884, 282.4978, 
    282.4072, 282.3167, 282.2261, 282.1355, 282.0449, 281.9543, 281.8638, 
    281.7732, 281.6826, 281.6943, 281.7544, 281.8145, 281.8745, 281.9346, 
    281.9946, 282.0547, 282.1147, 282.1748, 282.2349, 282.2949, 282.355, 
    282.415, 282.4844, 282.5732, 282.6643, 282.7581, 282.8542, 282.9531, 
    283.0547, 283.1592, 283.2668, 283.3777, 283.4917, 283.6091, 283.7302, 
    283.8542, 283.9014, 283.9548, 284.0156, 284.0854, 285.7424, 285.8472, 
    285.9377, 286.0171, 286.0869, 286.1492, 286.2046, 286.2546, 286.2998, 
    286.291, 286.2549, 286.2151, 286.1709, 286.1211, 286.0649, 286.0012, 
    285.928, 284.5112, 284.4478, 284.3931, 284.345, 284.3027, 284.2354, 
    284.1155, 283.9995, 283.887, 283.7776, 283.6714, 283.5684, 283.468, 
    283.3706, 283.2756, 283.1833, 283.0935, 283.0061, 282.9224, 282.936, 
    282.95, 282.9639, 282.9778, 282.9915, 283.0054, 283.0193, 283.0332, 
    283.0469, 283.0608, 283.0747, 283.0884, 283.1023, 283.0466, 282.958, 
    282.8696, 282.7812, 282.6926, 282.6042, 282.5159, 282.4272, 282.3389, 
    282.2505, 282.1619, 282.0735, 281.9851, 281.927, 281.9255, 281.9241, 
    281.9226, 281.9211, 281.9199, 281.9185, 281.917, 281.9155, 281.9143, 
    281.9128, 281.9114, 281.9099, 281.9092, 281.9436, 281.978, 282.0125, 
    282.0469, 282.0813, 282.1157, 282.1501, 282.1846, 282.2192, 282.2537, 
    282.2881, 282.3225, 282.3569, 282.3735, 282.3821, 282.3906, 282.3989, 
    282.4075, 282.416, 282.4243, 282.4329, 282.4414, 282.4497, 282.4583, 
    282.4668, 282.4751, 282.449, 282.3582, 282.2676, 282.1768, 282.0859, 
    281.9954, 281.9045, 281.8137, 281.7231, 281.6323, 281.5415, 281.4507, 
    281.3601, 281.2705, 281.2612, 281.2517, 281.2422, 281.2329, 281.2234, 
    281.2139, 281.2046, 281.1951, 281.1855, 281.1763, 281.1667, 281.1572, 
    281.1479, 281.1628, 281.1919, 281.2253, 281.2639, 281.3088, 282.4663, 
    282.5437, 282.6069, 282.6597, 282.7043, 282.7427, 282.7759, 282.8049, 
    282.8264, 282.8394, 282.8523, 282.8652, 282.8784, 282.8914, 282.9043, 
    282.9172, 282.9302, 282.9431, 282.9561, 282.969, 282.9819, 282.9939, 
    282.9502, 282.9065, 282.8628, 282.8191, 282.7751, 282.7314, 282.6877, 
    282.644, 282.6003, 282.5566, 282.5127, 282.469, 282.4253, 282.377, 
    282.321, 282.2571, 282.1833, 282.0972, 281.9954, 279.7285,
  280.0696, 280.2549, 280.4402, 280.6257, 280.811, 280.9966, 281.1819, 
    281.3672, 281.5527, 281.738, 281.9233, 282.1089, 282.2769, 282.4119, 
    282.5466, 282.6816, 282.8164, 282.9514, 283.0864, 283.2212, 283.3562, 
    283.4912, 283.626, 283.761, 283.8958, 284.0291, 284.0022, 283.9756, 
    283.949, 283.9224, 283.8958, 283.8689, 283.8423, 283.8157, 283.7891, 
    283.7625, 283.7356, 283.709, 283.6824, 283.7178, 283.7827, 283.8479, 
    283.9128, 283.9778, 284.0427, 284.1079, 284.1729, 284.2378, 284.3027, 
    284.3679, 284.4329, 284.4978, 284.5059, 284.406, 284.3062, 284.2063, 
    284.1064, 284.0066, 283.907, 283.8071, 283.7073, 283.6074, 283.5076, 
    283.4077, 283.3079, 283.208, 283.1047, 283.0017, 282.8987, 282.7957, 
    282.6926, 282.5894, 282.4863, 282.3833, 282.2803, 282.1772, 282.074, 
    281.9709, 281.8679, 281.8652, 281.9102, 281.9551, 281.9998, 282.0447, 
    282.0896, 282.1345, 282.1792, 282.2241, 282.269, 282.3137, 282.3586, 
    282.4036, 282.4609, 282.5449, 282.6323, 282.7241, 282.8201, 282.9207, 
    283.0264, 283.1375, 283.2542, 283.3774, 283.5073, 283.6445, 283.7898, 
    283.9424, 283.9988, 284.0618, 284.1331, 284.2139, 285.8608, 285.9629, 
    286.0544, 286.1372, 286.2122, 286.2805, 286.3433, 286.4006, 286.4539, 
    286.4434, 286.4019, 286.3567, 286.3076, 286.2537, 286.1946, 286.1292, 
    286.0569, 284.6345, 284.5608, 284.4963, 284.4395, 284.3889, 284.3083, 
    284.1682, 284.0359, 283.9109, 283.7925, 283.6804, 283.5737, 283.4724, 
    283.376, 283.2839, 283.1963, 283.1125, 283.0325, 282.9568, 282.9604, 
    282.9639, 282.9675, 282.9712, 282.9746, 282.9783, 282.9817, 282.9854, 
    282.9888, 282.9924, 282.9961, 282.9995, 283.0032, 282.9485, 282.8667, 
    282.7849, 282.7031, 282.6216, 282.5398, 282.458, 282.3762, 282.2944, 
    282.2126, 282.1309, 282.0491, 281.9673, 281.9146, 281.9158, 281.917, 
    281.9182, 281.9194, 281.9207, 281.9219, 281.9231, 281.9243, 281.9255, 
    281.9268, 281.928, 281.9292, 281.9312, 281.967, 282.0032, 282.0391, 
    282.0752, 282.1111, 282.1472, 282.1831, 282.2192, 282.2551, 282.2913, 
    282.3271, 282.3633, 282.3992, 282.4126, 282.4153, 282.418, 282.4207, 
    282.4233, 282.4263, 282.429, 282.4316, 282.4343, 282.437, 282.4397, 
    282.4426, 282.4453, 282.4182, 282.3354, 282.2527, 282.1699, 282.0872, 
    282.0044, 281.9216, 281.8389, 281.7561, 281.6733, 281.5906, 281.5078, 
    281.425, 281.3435, 281.335, 281.3267, 281.3181, 281.3098, 281.3013, 
    281.293, 281.2844, 281.2761, 281.2676, 281.2593, 281.2507, 281.2424, 
    281.2339, 281.2488, 281.2771, 281.3093, 281.3467, 281.3904, 282.5137, 
    282.5889, 282.6501, 282.7014, 282.7449, 282.782, 282.8142, 282.8423, 
    282.864, 282.8792, 282.894, 282.9089, 282.9238, 282.9387, 282.9539, 
    282.9688, 282.9836, 282.9985, 283.0134, 283.0286, 283.0435, 283.0574, 
    283.0151, 282.9731, 282.9309, 282.8887, 282.8467, 282.8044, 282.7622, 
    282.72, 282.678, 282.6357, 282.5935, 282.5515, 282.5093, 282.4607, 
    282.4031, 282.3374, 282.2615, 282.1729, 282.0684, 279.7388,
  280.1682, 280.3521, 280.5359, 280.72, 280.9038, 281.0876, 281.2717, 
    281.4556, 281.6394, 281.8235, 282.0073, 282.1912, 282.3564, 282.4863, 
    282.6162, 282.7458, 282.8757, 283.0054, 283.1353, 283.2651, 283.3948, 
    283.5247, 283.6543, 283.7842, 283.9141, 284.042, 284.0122, 283.9824, 
    283.9526, 283.9229, 283.8931, 283.863, 283.8333, 283.8035, 283.7737, 
    283.7439, 283.7141, 283.6843, 283.6545, 283.6821, 283.7373, 283.7922, 
    283.8474, 283.9026, 283.9575, 284.0127, 284.0676, 284.1228, 284.178, 
    284.2329, 284.2881, 284.343, 284.3579, 284.2964, 284.2346, 284.1729, 
    284.1113, 284.0496, 283.988, 283.9263, 283.8647, 283.803, 283.7412, 
    283.6797, 283.6179, 283.5557, 283.4402, 283.3245, 283.209, 283.0933, 
    282.9778, 282.8623, 282.7466, 282.6311, 282.5154, 282.3999, 282.2842, 
    282.1687, 282.0532, 282.0361, 282.0659, 282.0955, 282.1252, 282.1548, 
    282.1843, 282.2141, 282.2437, 282.2734, 282.303, 282.3328, 282.3623, 
    282.3921, 282.4375, 282.5156, 282.5991, 282.688, 282.783, 282.8848, 
    282.9941, 283.1121, 283.2393, 283.377, 283.5269, 283.6902, 283.8694, 
    284.0645, 284.1318, 284.207, 284.2908, 284.3853, 285.957, 286.0601, 
    286.1555, 286.2441, 286.3267, 286.4038, 286.4758, 286.5435, 286.6069, 
    286.5942, 286.5444, 286.4912, 286.4346, 286.374, 286.3088, 286.239, 
    286.1636, 284.7979, 284.7119, 284.636, 284.5681, 284.5076, 284.408, 
    284.2375, 284.0825, 283.9407, 283.8105, 283.6907, 283.5801, 283.4773, 
    283.3818, 283.293, 283.21, 283.1321, 283.0591, 282.9915, 282.9846, 
    282.978, 282.9712, 282.9646, 282.9578, 282.9509, 282.9443, 282.9375, 
    282.9309, 282.9241, 282.9172, 282.9106, 282.9038, 282.8506, 282.7754, 
    282.7004, 282.6252, 282.5503, 282.4751, 282.4001, 282.325, 282.25, 
    282.1748, 282.0999, 282.0247, 281.9497, 281.9021, 281.906, 281.9099, 
    281.9138, 281.9177, 281.9214, 281.9253, 281.9292, 281.9331, 281.937, 
    281.9409, 281.9448, 281.9487, 281.9531, 281.9907, 282.0283, 282.0657, 
    282.1033, 282.1409, 282.1785, 282.2161, 282.2537, 282.2913, 282.3289, 
    282.3665, 282.4041, 282.4414, 282.4514, 282.4485, 282.4453, 282.4424, 
    282.4395, 282.4363, 282.4333, 282.4304, 282.4275, 282.4243, 282.4214, 
    282.4185, 282.4153, 282.3872, 282.3125, 282.2378, 282.1631, 282.0881, 
    282.0134, 281.9387, 281.8638, 281.7891, 281.7144, 281.6394, 281.5647, 
    281.49, 281.4163, 281.4089, 281.4014, 281.394, 281.3867, 281.3792, 
    281.3718, 281.3645, 281.3572, 281.3496, 281.3423, 281.335, 281.3274, 
    281.3201, 281.3347, 281.3621, 281.3936, 281.4297, 281.4719, 282.561, 
    282.634, 282.6936, 282.7432, 282.7852, 282.8213, 282.8525, 282.8799, 
    282.9019, 282.9187, 282.9355, 282.9526, 282.9695, 282.9863, 283.0032, 
    283.0203, 283.0371, 283.054, 283.071, 283.0879, 283.1047, 283.1208, 
    283.0801, 283.0396, 282.999, 282.9585, 282.918, 282.8772, 282.8367, 
    282.7961, 282.7556, 282.7151, 282.6743, 282.6338, 282.5933, 282.5442, 
    282.4851, 282.4175, 282.3396, 282.2488, 282.1411, 279.7493,
  280.2668, 280.4492, 280.6316, 280.8142, 280.9966, 281.179, 281.3613, 
    281.5439, 281.7263, 281.9087, 282.0913, 282.2737, 282.4363, 282.5608, 
    282.6855, 282.8101, 282.9348, 283.0596, 283.1841, 283.3088, 283.4333, 
    283.5581, 283.6829, 283.8074, 283.9321, 284.0549, 284.022, 283.989, 
    283.9561, 283.9231, 283.8901, 283.8572, 283.8242, 283.7913, 283.7583, 
    283.7253, 283.6924, 283.6594, 283.6265, 283.6465, 283.6917, 283.7368, 
    283.782, 283.8271, 283.8723, 283.9175, 283.9626, 284.0078, 284.053, 
    284.0981, 284.1433, 284.1885, 284.21, 284.1865, 284.1631, 284.1394, 
    284.116, 284.0925, 284.0691, 284.0457, 284.022, 283.9985, 283.9751, 
    283.9517, 283.9282, 283.9033, 283.7754, 283.6472, 283.5193, 283.3911, 
    283.2629, 283.135, 283.0068, 282.8787, 282.7507, 282.6226, 282.4944, 
    282.3665, 282.2383, 282.207, 282.2214, 282.2358, 282.2505, 282.2649, 
    282.2793, 282.2937, 282.3083, 282.3228, 282.3372, 282.3516, 282.3662, 
    282.3806, 282.4138, 282.4858, 282.5642, 282.6494, 282.7427, 282.8447, 
    282.9573, 283.082, 283.2209, 283.3765, 285.1809, 285.2654, 285.3406, 
    285.4084, 285.5488, 285.6812, 285.8062, 285.9243, 286.0366, 286.1428, 
    286.2441, 286.3403, 286.4319, 286.5193, 286.6028, 286.6826, 286.759, 
    286.7432, 286.6826, 286.6191, 286.553, 286.4834, 286.4106, 286.3342, 
    286.2537, 286.1689, 286.0798, 285.9856, 285.886, 285.7805, 285.6882, 
    285.6262, 285.5566, 285.478, 285.3882, 285.2847, 285.1641, 285.022, 
    284.8518, 284.6448, 284.387, 284.0574, 283.0864, 283.0261, 283.009, 
    282.9919, 282.9749, 282.958, 282.9409, 282.9238, 282.9067, 282.8896, 
    282.8728, 282.8557, 282.8386, 282.8215, 282.8047, 282.7527, 282.6841, 
    282.6157, 282.5474, 282.479, 282.4106, 282.3423, 282.2739, 282.2056, 
    282.1372, 282.0688, 282.0002, 281.9319, 281.8896, 281.8962, 281.9028, 
    281.9092, 281.9158, 281.9224, 281.929, 281.9353, 281.9419, 281.9485, 
    281.9548, 281.9614, 281.968, 281.9751, 282.0142, 282.0532, 282.0925, 
    282.1316, 282.1707, 282.21, 282.249, 282.2881, 282.3271, 282.3665, 
    282.4055, 282.4446, 282.4839, 282.4902, 282.4817, 282.4729, 282.4641, 
    282.4553, 282.4465, 282.438, 282.4292, 282.4204, 282.4116, 282.4028, 
    282.3943, 282.3855, 282.3564, 282.2898, 282.2229, 282.156, 282.0894, 
    282.0225, 281.9558, 281.8889, 281.822, 281.7554, 281.6885, 281.6216, 
    281.5549, 281.489, 281.4827, 281.4763, 281.47, 281.4636, 281.4573, 
    281.4509, 281.4443, 281.438, 281.4316, 281.4253, 281.4189, 281.4126, 
    281.4062, 281.4204, 281.447, 281.4775, 281.5125, 281.5535, 282.6086, 
    282.6792, 282.7368, 282.7849, 282.8257, 282.8606, 282.8909, 282.9172, 
    282.9395, 282.9583, 282.9773, 282.9961, 283.0151, 283.0339, 283.0527, 
    283.0718, 283.0906, 283.1096, 283.1284, 283.1472, 283.1663, 283.1841, 
    283.1453, 283.1062, 283.0671, 283.0281, 282.9893, 282.9502, 282.9111, 
    282.8723, 282.8333, 282.7942, 282.7551, 282.7163, 282.6772, 282.6277, 
    282.5671, 282.4978, 282.4177, 282.3245, 282.2141, 279.7595,
  280.3655, 280.5464, 280.7273, 280.9084, 281.0894, 281.2703, 281.4512, 
    281.6321, 281.8132, 281.9941, 282.175, 282.356, 282.5159, 282.6353, 
    282.7549, 282.8745, 282.9939, 283.1135, 283.2332, 283.3525, 283.4722, 
    283.5916, 283.7112, 283.8308, 283.9502, 284.0681, 284.032, 283.9958, 
    283.9597, 283.9236, 283.8875, 283.8513, 283.8154, 283.7793, 283.7432, 
    283.707, 283.6709, 283.6348, 283.5986, 283.6108, 283.6462, 283.6814, 
    283.7166, 283.752, 283.7871, 283.8223, 283.8577, 283.8928, 283.928, 
    283.9634, 283.9985, 284.0337, 284.062, 284.0767, 284.0913, 284.106, 
    284.1208, 284.1355, 284.1501, 284.1648, 284.1794, 284.1943, 284.209, 
    284.2236, 284.2383, 284.2512, 284.1106, 283.97, 283.8293, 283.6887, 
    283.5483, 283.4077, 283.2671, 283.1265, 282.9858, 282.8452, 282.7046, 
    282.5642, 282.4236, 282.3779, 282.3772, 282.3765, 282.3757, 282.375, 
    282.3743, 282.3735, 282.3728, 282.3721, 282.3713, 282.3706, 282.3699, 
    282.3691, 282.3899, 282.4553, 282.5278, 282.6084, 282.6985, 282.7998, 
    282.915, 283.0466, 283.1985, 283.376, 285.291, 285.3679, 285.4355, 
    285.4966, 285.6252, 285.7502, 285.8716, 285.989, 286.1033, 286.2144, 
    286.3223, 286.427, 286.5291, 286.6282, 286.7249, 286.8188, 286.9104, 
    286.8904, 286.8167, 286.7412, 286.6636, 286.5837, 286.5017, 286.4175, 
    286.3306, 286.2415, 286.1494, 286.0549, 285.9573, 285.8567, 285.772, 
    285.7173, 285.6555, 285.585, 285.5039, 285.4094, 285.2983, 285.1653, 
    285.0037, 284.8025, 284.5461, 284.207, 283.1143, 283.0605, 283.0332, 
    283.0059, 282.9788, 282.9514, 282.9241, 282.8967, 282.8694, 282.842, 
    282.8147, 282.7874, 282.76, 282.7327, 282.7053, 282.6545, 282.5928, 
    282.5312, 282.4695, 282.4077, 282.3462, 282.2844, 282.2227, 282.1611, 
    282.0994, 282.0376, 281.9761, 281.9143, 281.8772, 281.8865, 281.8955, 
    281.9048, 281.9141, 281.9231, 281.9324, 281.9414, 281.9507, 281.9597, 
    281.969, 281.9783, 281.9873, 281.9971, 282.0376, 282.0784, 282.1191, 
    282.1599, 282.2004, 282.2412, 282.282, 282.3225, 282.3633, 282.4041, 
    282.4448, 282.4854, 282.5261, 282.5293, 282.5146, 282.5002, 282.4858, 
    282.4714, 282.4568, 282.4424, 282.428, 282.4136, 282.3989, 282.3845, 
    282.3701, 282.3555, 282.3257, 282.2668, 282.208, 282.1492, 282.0903, 
    282.0315, 281.9727, 281.9138, 281.8552, 281.7964, 281.7375, 281.6787, 
    281.6199, 281.562, 281.5566, 281.5513, 281.5459, 281.5405, 281.5352, 
    281.5298, 281.5244, 281.519, 281.5137, 281.5083, 281.5029, 281.4976, 
    281.4922, 281.5063, 281.5322, 281.5615, 281.5955, 281.635, 282.656, 
    282.7244, 282.78, 282.8267, 282.866, 282.8999, 282.9292, 282.9548, 
    282.9771, 282.998, 283.0188, 283.0398, 283.0605, 283.0815, 283.1023, 
    283.1233, 283.144, 283.165, 283.1858, 283.2068, 283.2275, 283.2476, 
    283.2102, 283.1726, 283.1353, 283.0979, 283.0605, 283.0232, 282.9856, 
    282.9482, 282.9109, 282.8735, 282.8359, 282.7986, 282.7612, 282.7112, 
    282.6489, 282.5779, 282.4958, 282.4001, 282.2871, 279.7698,
  280.4641, 280.6436, 280.8232, 281.0027, 281.1821, 281.3616, 281.541, 
    281.7205, 281.8999, 282.0793, 282.259, 282.4385, 282.5955, 282.71, 
    282.8242, 282.9387, 283.0532, 283.1675, 283.282, 283.3962, 283.5107, 
    283.6252, 283.7395, 283.854, 283.9683, 284.0811, 284.0417, 284.0027, 
    283.9634, 283.9241, 283.8848, 283.8455, 283.8064, 283.7671, 283.7278, 
    283.6885, 283.6494, 283.6101, 283.5708, 283.5754, 283.6006, 283.626, 
    283.6514, 283.6765, 283.7019, 283.7273, 283.7524, 283.7778, 283.8032, 
    283.8284, 283.8538, 283.8792, 283.9138, 283.9668, 284.0198, 284.0725, 
    284.1255, 284.1785, 284.2312, 284.2842, 284.3369, 284.3899, 284.4429, 
    284.4956, 284.5486, 284.5989, 284.4458, 284.2927, 284.1396, 283.9866, 
    283.8335, 283.6804, 283.5273, 283.3743, 283.2212, 283.0679, 282.9148, 
    282.7617, 282.6086, 282.5488, 282.5327, 282.5168, 282.501, 282.4851, 
    282.4692, 282.4531, 282.4373, 282.4214, 282.4055, 282.3896, 282.3735, 
    282.3577, 282.366, 282.4241, 282.4897, 282.5645, 282.6501, 282.7493, 
    282.8652, 283.0034, 283.1702, 283.3752, 285.376, 285.4465, 285.5081, 
    285.5632, 285.6848, 285.8054, 285.9248, 286.0432, 286.1604, 286.2764, 
    286.3916, 286.5056, 286.6187, 286.7307, 286.8418, 286.9519, 287.061, 
    287.0356, 286.947, 286.8574, 286.7668, 286.6758, 286.5837, 286.491, 
    286.3972, 286.3027, 286.2073, 286.1108, 286.0137, 285.9155, 285.8354, 
    285.7869, 285.7314, 285.668, 285.5942, 285.5081, 285.4053, 285.2812, 
    285.1282, 284.9348, 284.6829, 284.3403, 283.1423, 283.0952, 283.0576, 
    283.02, 282.9824, 282.9448, 282.907, 282.8694, 282.8318, 282.7942, 
    282.7566, 282.719, 282.6814, 282.6438, 282.606, 282.5566, 282.5017, 
    282.4465, 282.3916, 282.3367, 282.2815, 282.2266, 282.1716, 282.1167, 
    282.0615, 282.0066, 281.9517, 281.8965, 281.8647, 281.8767, 281.8884, 
    281.9004, 281.9121, 281.9238, 281.9358, 281.9475, 281.9595, 281.9712, 
    281.9832, 281.9949, 282.0066, 282.019, 282.0613, 282.1035, 282.1458, 
    282.188, 282.2302, 282.2725, 282.3149, 282.3572, 282.3994, 282.4417, 
    282.4839, 282.5261, 282.5684, 282.5681, 282.5479, 282.5276, 282.5076, 
    282.4873, 282.467, 282.4468, 282.4268, 282.4065, 282.3862, 282.366, 
    282.3459, 282.3257, 282.2949, 282.2439, 282.1931, 282.1423, 282.0916, 
    282.0405, 281.9897, 281.939, 281.8882, 281.8374, 281.7864, 281.7356, 
    281.6848, 281.6348, 281.6304, 281.626, 281.6218, 281.6174, 281.613, 
    281.6086, 281.6045, 281.6001, 281.5957, 281.5913, 281.5872, 281.5828, 
    281.5784, 281.5923, 281.6172, 281.6455, 281.6785, 281.7168, 282.7034, 
    282.7695, 282.8235, 282.8684, 282.9065, 282.9392, 282.9675, 282.9922, 
    283.0146, 283.0376, 283.0605, 283.0833, 283.1062, 283.1292, 283.1519, 
    283.1748, 283.1975, 283.2205, 283.2434, 283.2661, 283.2891, 283.3108, 
    283.2751, 283.2393, 283.2034, 283.1677, 283.1318, 283.0959, 283.0601, 
    283.0244, 282.9885, 282.9526, 282.9167, 282.8811, 282.8452, 282.7947, 
    282.731, 282.6582, 282.5742, 282.4761, 282.3601, 279.78,
  280.6221, 280.8015, 280.9812, 281.1609, 281.3403, 281.52, 281.6997, 
    281.8792, 282.0588, 282.2385, 282.418, 282.5977, 282.7524, 282.8596, 
    282.967, 283.0742, 283.1816, 283.2888, 283.3962, 283.5034, 283.6108, 
    283.718, 283.8254, 283.9326, 284.04, 284.1458, 284.1033, 284.0605, 
    284.0181, 283.9756, 283.9331, 283.8904, 283.8479, 283.8054, 283.7629, 
    283.7202, 283.6777, 283.6353, 283.5928, 283.5913, 283.6094, 283.6274, 
    283.6455, 283.6636, 283.6816, 283.6997, 283.7178, 283.7358, 283.7539, 
    283.772, 283.79, 283.8081, 283.8447, 283.9167, 283.9895, 284.0627, 
    284.1365, 284.2109, 284.2861, 284.3621, 284.4385, 284.5154, 284.5933, 
    284.6716, 284.7507, 284.8276, 284.6687, 284.5098, 284.3508, 284.1919, 
    284.033, 283.874, 283.7153, 283.5564, 283.3975, 283.2385, 283.0796, 
    282.9207, 282.7617, 282.6948, 282.6714, 282.6479, 282.6245, 282.6013, 
    282.5779, 282.5544, 282.531, 282.5078, 282.4844, 282.4609, 282.4377, 
    282.4143, 282.4175, 282.4756, 282.5417, 282.6174, 282.7053, 282.8083, 
    282.9309, 283.0791, 283.262, 283.4929, 285.5461, 285.603, 285.6533, 
    285.6987, 285.8096, 285.9202, 286.031, 286.1416, 286.2524, 286.3633, 
    286.4739, 286.5847, 286.6953, 286.8062, 286.917, 287.0276, 287.1384, 
    287.1101, 287.0166, 286.9231, 286.8296, 286.7361, 286.6426, 286.5491, 
    286.4556, 286.3618, 286.2683, 286.1748, 286.0813, 285.9878, 285.9121, 
    285.8657, 285.8132, 285.7527, 285.6824, 285.5996, 285.5007, 285.3806, 
    285.2317, 285.0422, 284.7925, 284.4492, 283.1995, 283.1553, 283.1047, 
    283.0542, 283.0037, 282.9531, 282.9026, 282.8518, 282.8013, 282.7507, 
    282.7002, 282.6497, 282.5991, 282.5486, 282.4978, 282.4502, 282.4041, 
    282.3577, 282.3113, 282.2651, 282.2188, 282.1724, 282.1262, 282.0798, 
    282.0334, 281.9873, 281.9409, 281.8945, 281.8687, 281.8809, 281.8933, 
    281.9055, 281.918, 281.9302, 281.9424, 281.9548, 281.967, 281.9795, 
    281.9917, 282.0039, 282.0164, 282.0291, 282.0693, 282.1096, 282.1497, 
    282.1899, 282.2302, 282.2705, 282.3108, 282.3511, 282.3911, 282.4314, 
    282.4717, 282.512, 282.5522, 282.552, 282.5332, 282.5144, 282.4954, 
    282.4766, 282.4578, 282.4387, 282.4199, 282.4011, 282.3821, 282.3633, 
    282.3445, 282.3254, 282.2979, 282.2539, 282.2095, 282.1646, 282.1194, 
    282.074, 282.0281, 281.9817, 281.9348, 281.8877, 281.8403, 281.7922, 
    281.7439, 281.6958, 281.6921, 281.6882, 281.6846, 281.6807, 281.677, 
    281.6733, 281.6694, 281.6658, 281.6619, 281.6582, 281.6545, 281.6506, 
    281.647, 281.6616, 281.6873, 281.7168, 281.7507, 281.79, 282.7991, 
    282.8511, 282.8948, 282.9316, 282.9636, 282.9912, 283.0154, 283.0369, 
    283.0576, 283.0806, 283.1035, 283.1265, 283.1494, 283.1724, 283.1953, 
    283.2183, 283.2412, 283.2642, 283.2871, 283.3101, 283.333, 283.355, 
    283.3208, 283.2869, 283.2527, 283.2185, 283.1843, 283.1504, 283.1162, 
    283.082, 283.0479, 283.0137, 282.9797, 282.9456, 282.9114, 282.8611, 
    282.7966, 282.7229, 282.6377, 282.5386, 282.4211, 279.8105,
  280.8423, 281.0239, 281.2053, 281.3867, 281.5681, 281.7495, 281.9309, 
    282.1125, 282.2939, 282.4753, 282.6567, 282.8381, 282.991, 283.0891, 
    283.1873, 283.2854, 283.3835, 283.4814, 283.5796, 283.6777, 283.7759, 
    283.874, 283.9722, 284.0703, 284.1685, 284.2649, 284.219, 284.1729, 
    284.127, 284.0811, 284.0349, 283.989, 283.9431, 283.897, 283.8511, 
    283.8052, 283.759, 283.7131, 283.6672, 283.6616, 283.6753, 283.689, 
    283.7026, 283.7163, 283.73, 283.7437, 283.7573, 283.771, 283.7847, 
    283.7983, 283.812, 283.8257, 283.8589, 283.9302, 284.0032, 284.0784, 
    284.1553, 284.2344, 284.3159, 284.3994, 284.4854, 284.5737, 284.6648, 
    284.7585, 284.8552, 284.9517, 284.7942, 284.6367, 284.4792, 284.3218, 
    284.1643, 284.0068, 283.8494, 283.6919, 283.5344, 283.377, 283.2195, 
    283.062, 282.9045, 282.8389, 282.8164, 282.7939, 282.7712, 282.7488, 
    282.7263, 282.7039, 282.6814, 282.6589, 282.6365, 282.614, 282.5916, 
    282.5688, 282.5757, 282.6428, 282.7188, 282.8052, 282.905, 283.021, 
    283.1577, 283.321, 283.52, 283.7676, 285.8091, 285.8491, 285.8853, 
    285.9189, 286.0127, 286.1067, 286.2004, 286.2942, 286.3882, 286.4819, 
    286.5759, 286.6697, 286.7637, 286.8574, 286.9514, 287.0452, 287.1392, 
    287.1108, 287.0254, 286.9397, 286.8542, 286.7688, 286.6831, 286.5977, 
    286.512, 286.4265, 286.3411, 286.2554, 286.1699, 286.0842, 286.0137, 
    285.9673, 285.9143, 285.8535, 285.7827, 285.6995, 285.6001, 285.4795, 
    285.3298, 285.1392, 284.8884, 284.5432, 283.2871, 283.2424, 283.176, 
    283.1099, 283.0435, 282.9771, 282.9109, 282.8445, 282.7783, 282.7119, 
    282.6455, 282.5793, 282.5129, 282.4468, 282.3804, 282.335, 282.2996, 
    282.2642, 282.2285, 282.1931, 282.1577, 282.1221, 282.0867, 282.0513, 
    282.0156, 281.9802, 281.9446, 281.9092, 281.8896, 281.9001, 281.9106, 
    281.9211, 281.9316, 281.9421, 281.9526, 281.9631, 281.9736, 281.9841, 
    281.9946, 282.0051, 282.0156, 282.0264, 282.0608, 282.0952, 282.1296, 
    282.1641, 282.1985, 282.2329, 282.2673, 282.3018, 282.3362, 282.3706, 
    282.405, 282.4395, 282.4739, 282.478, 282.468, 282.4578, 282.4478, 
    282.4375, 282.4275, 282.4175, 282.4072, 282.3972, 282.387, 282.377, 
    282.3669, 282.3567, 282.3372, 282.2993, 282.2603, 282.2205, 282.1792, 
    282.1372, 282.0938, 282.0493, 282.0037, 281.9565, 281.908, 281.8582, 
    281.8066, 281.7544, 281.7507, 281.7471, 281.7434, 281.7397, 281.7361, 
    281.7324, 281.729, 281.7253, 281.7217, 281.718, 281.7144, 281.7107, 
    281.707, 281.7236, 281.7527, 281.7854, 281.823, 281.8665, 282.9233, 
    282.9568, 282.9858, 283.0115, 283.0339, 283.0542, 283.0723, 283.0886, 
    283.1057, 283.127, 283.1479, 283.1689, 283.1899, 283.2112, 283.2322, 
    283.2532, 283.2742, 283.2954, 283.3164, 283.3374, 283.3584, 283.3787, 
    283.3464, 283.314, 283.2817, 283.2495, 283.2173, 283.1848, 283.1526, 
    283.1204, 283.0881, 283.0557, 283.0234, 282.9912, 282.959, 282.9092, 
    282.8447, 282.7712, 282.6863, 282.5872, 282.47, 279.8621,
  281.0627, 281.2461, 281.4292, 281.6125, 281.7959, 281.9792, 282.1624, 
    282.3457, 282.5291, 282.7122, 282.8955, 283.0789, 283.2295, 283.3186, 
    283.4075, 283.4963, 283.5852, 283.6743, 283.7632, 283.8521, 283.9409, 
    284.0298, 284.1189, 284.2078, 284.2966, 284.384, 284.3347, 284.2852, 
    284.2358, 284.1863, 284.137, 284.0876, 284.0381, 283.9888, 283.9392, 
    283.8899, 283.8403, 283.791, 283.7417, 283.7319, 283.7412, 283.7505, 
    283.7598, 283.769, 283.7783, 283.7876, 283.7969, 283.8062, 283.8154, 
    283.8247, 283.834, 283.8433, 283.873, 283.9438, 284.0176, 284.0947, 
    284.1755, 284.2603, 284.3491, 284.4424, 284.5405, 284.6438, 284.7527, 
    284.8677, 284.9895, 285.1147, 284.9592, 284.8037, 284.6482, 284.4927, 
    284.3372, 284.1816, 284.0261, 283.8706, 283.7151, 283.5596, 283.4041, 
    283.2485, 283.093, 283.0286, 283.0073, 282.9858, 282.9646, 282.9434, 
    282.9221, 282.9006, 282.8794, 282.8582, 282.8367, 282.8154, 282.7942, 
    282.7727, 282.7837, 282.8616, 282.9487, 283.0476, 283.1604, 283.2905, 
    283.4419, 283.6204, 283.8342, 284.0947, 286.0566, 286.0862, 286.1133, 
    286.1389, 286.2161, 286.293, 286.3699, 286.447, 286.5239, 286.6008, 
    286.678, 286.7549, 286.8318, 286.9087, 286.9858, 287.0627, 287.1396, 
    287.1116, 287.0339, 286.9565, 286.8789, 286.8013, 286.7239, 286.6462, 
    286.5686, 286.491, 286.4136, 286.3359, 286.2583, 286.1807, 286.1152, 
    286.0686, 286.0154, 285.9543, 285.8831, 285.7996, 285.6997, 285.5784, 
    285.428, 285.2363, 284.9841, 284.6372, 283.3745, 283.3293, 283.2473, 
    283.1653, 283.0833, 283.0012, 282.9192, 282.8372, 282.7551, 282.6731, 
    282.5911, 282.509, 282.427, 282.345, 282.2629, 282.22, 282.1953, 
    282.1707, 282.146, 282.1211, 282.0964, 282.0718, 282.0471, 282.0225, 
    281.9978, 281.9731, 281.9485, 281.9238, 281.9106, 281.9194, 281.9282, 
    281.9368, 281.9456, 281.9541, 281.9629, 281.9714, 281.9802, 281.9888, 
    281.9976, 282.0061, 282.0149, 282.0239, 282.0525, 282.0811, 282.1096, 
    282.1382, 282.167, 282.1956, 282.2241, 282.2527, 282.2812, 282.3101, 
    282.3386, 282.3672, 282.3958, 282.4041, 282.4026, 282.4014, 282.3999, 
    282.3987, 282.3972, 282.396, 282.3948, 282.3933, 282.3921, 282.3906, 
    282.3894, 282.3879, 282.3767, 282.3457, 282.3132, 282.2795, 282.2441, 
    282.207, 282.168, 282.1272, 282.084, 282.0388, 281.991, 281.9407, 
    281.8872, 281.8318, 281.8281, 281.8247, 281.8213, 281.8176, 281.8142, 
    281.8108, 281.8071, 281.8037, 281.8, 281.7966, 281.7932, 281.7896, 
    281.7861, 281.8052, 281.8379, 281.8745, 281.916, 281.9639, 283.0247, 
    283.0461, 283.0657, 283.0833, 283.0994, 283.114, 283.1274, 283.1399, 
    283.1541, 283.1731, 283.1924, 283.2114, 283.2307, 283.2498, 283.269, 
    283.2881, 283.3074, 283.3264, 283.3457, 283.3647, 283.384, 283.4023, 
    283.3718, 283.3413, 283.311, 283.2805, 283.25, 283.2195, 283.1892, 
    283.1587, 283.1282, 283.0977, 283.0674, 283.0369, 283.0063, 282.9573, 
    282.8928, 282.8193, 282.7346, 282.6355, 282.5186, 279.9136,
  281.2832, 281.4683, 281.6533, 281.8384, 282.0237, 282.2087, 282.3938, 
    282.5789, 282.7639, 282.9492, 283.1343, 283.3193, 283.4683, 283.5479, 
    283.6277, 283.7073, 283.7871, 283.8669, 283.9465, 284.0264, 284.106, 
    284.1858, 284.2654, 284.3452, 284.425, 284.5032, 284.4504, 284.3975, 
    284.3447, 284.2917, 284.239, 284.186, 284.1333, 284.0803, 284.0276, 
    283.9746, 283.9219, 283.8689, 283.8162, 283.8022, 283.8071, 283.812, 
    283.8169, 283.8218, 283.8267, 283.8318, 283.8367, 283.8416, 283.8464, 
    283.8513, 283.8562, 283.8611, 283.8875, 283.9578, 284.0327, 284.1125, 
    284.1978, 284.2891, 284.387, 284.4924, 284.6062, 284.7292, 284.863, 
    285.0088, 285.1685, 285.3396, 285.1868, 285.0339, 284.8811, 284.728, 
    284.5752, 284.4224, 284.2695, 284.1167, 283.9639, 283.811, 283.6582, 
    283.5054, 283.3525, 283.29, 283.2703, 283.2505, 283.231, 283.2112, 
    283.1914, 283.1719, 283.1521, 283.1323, 283.1125, 283.093, 283.0732, 
    283.0535, 283.0696, 283.1597, 283.26, 283.3723, 283.499, 283.6433, 
    283.8086, 284, 284.2246, 284.4915, 286.2905, 286.3147, 286.3374, 
    286.3591, 286.4192, 286.4792, 286.5396, 286.5996, 286.6597, 286.7197, 
    286.7798, 286.8398, 286.9001, 286.9602, 287.0203, 287.0803, 287.1404, 
    287.1123, 287.0427, 286.9731, 286.9036, 286.834, 286.7644, 286.6948, 
    286.6252, 286.5557, 286.4861, 286.4165, 286.3469, 286.2773, 286.2168, 
    286.1699, 286.1165, 286.0549, 285.9836, 285.8994, 285.7991, 285.6772, 
    285.5259, 285.3335, 285.0798, 284.7312, 283.4619, 283.4165, 283.3186, 
    283.2209, 283.123, 283.0254, 282.9275, 282.8298, 282.7319, 282.6343, 
    282.5364, 282.4387, 282.3408, 282.2432, 282.1453, 282.1047, 282.0908, 
    282.0769, 282.0632, 282.0493, 282.0354, 282.0215, 282.0078, 281.9939, 
    281.98, 281.9661, 281.9524, 281.9385, 281.9319, 281.9387, 281.9456, 
    281.9524, 281.9592, 281.9661, 281.9729, 281.9797, 281.9868, 281.9937, 
    282.0005, 282.0073, 282.0142, 282.0212, 282.0439, 282.0669, 282.0896, 
    282.1125, 282.1353, 282.158, 282.1809, 282.2036, 282.2263, 282.2493, 
    282.272, 282.2949, 282.3176, 282.3298, 282.3374, 282.3447, 282.3523, 
    282.3596, 282.3672, 282.3745, 282.3821, 282.3894, 282.397, 282.4043, 
    282.4119, 282.4192, 282.4163, 282.3933, 282.3687, 282.3423, 282.3142, 
    282.2842, 282.252, 282.2173, 282.1799, 282.1394, 282.0952, 282.0474, 
    281.9949, 281.938, 281.9348, 281.9314, 281.9282, 281.9248, 281.9216, 
    281.9182, 281.915, 281.9116, 281.9084, 281.905, 281.9019, 281.8984, 
    281.8953, 281.917, 281.9536, 281.9944, 282.0403, 282.0923, 283.1086, 
    283.123, 283.1362, 283.1487, 283.1602, 283.1709, 283.1809, 283.1904, 
    283.2021, 283.2195, 283.2368, 283.2542, 283.2712, 283.2886, 283.3059, 
    283.3232, 283.3403, 283.3577, 283.375, 283.3921, 283.4094, 283.426, 
    283.3972, 283.3687, 283.3401, 283.3115, 283.283, 283.2542, 283.2256, 
    283.197, 283.1685, 283.1396, 283.1111, 283.0825, 283.054, 283.0054, 
    282.9412, 282.8677, 282.783, 282.6841, 282.5671, 279.9651,
  281.5034, 281.6904, 281.8774, 282.0645, 282.2512, 282.4382, 282.6252, 
    282.812, 282.999, 283.186, 283.373, 283.5598, 283.7068, 283.7773, 
    283.8479, 283.9185, 283.989, 284.0596, 284.1301, 284.2007, 284.271, 
    284.3416, 284.4121, 284.4827, 284.5532, 284.6223, 284.5662, 284.5098, 
    284.4536, 284.3972, 284.3408, 284.2847, 284.2283, 284.1721, 284.1157, 
    284.0593, 284.0032, 283.9468, 283.8906, 283.8728, 283.8733, 283.8738, 
    283.8743, 283.8748, 283.8752, 283.8757, 283.8762, 283.8767, 283.8772, 
    283.8777, 283.8782, 283.8787, 283.9019, 283.9722, 284.0483, 284.1311, 
    284.2217, 284.3208, 284.4302, 284.551, 284.6855, 284.8359, 285.0056, 
    285.1982, 285.4189, 285.6689, 285.52, 285.3711, 285.2219, 285.073, 
    284.9241, 284.7751, 284.6262, 284.4773, 284.3284, 284.1794, 284.0305, 
    283.8816, 283.7327, 283.6731, 283.6558, 283.6384, 283.6211, 283.6035, 
    283.5862, 283.5688, 283.5515, 283.5342, 283.5168, 283.4995, 283.4822, 
    283.4648, 283.4871, 283.5906, 283.7043, 283.8298, 283.9692, 284.1248, 
    284.2996, 284.4973, 284.7229, 284.9827, 286.5115, 286.5349, 286.5574, 
    286.5793, 286.6226, 286.6658, 286.709, 286.7522, 286.7954, 286.8386, 
    286.8818, 286.925, 286.9683, 287.0115, 287.0547, 287.0979, 287.1411, 
    287.113, 287.0515, 286.9897, 286.9282, 286.8667, 286.8049, 286.7434, 
    286.6819, 286.6201, 286.5586, 286.4971, 286.4353, 286.3738, 286.3186, 
    286.2715, 286.2175, 286.1558, 286.084, 285.9995, 285.8987, 285.7761, 
    285.624, 285.4304, 285.1758, 284.8252, 283.5496, 283.5034, 283.3899, 
    283.2764, 283.1628, 283.0493, 282.9358, 282.8225, 282.709, 282.5955, 
    282.4819, 282.3684, 282.2549, 282.1414, 282.0278, 281.9895, 281.9866, 
    281.9834, 281.9805, 281.9773, 281.9744, 281.9712, 281.9683, 281.9653, 
    281.9622, 281.9592, 281.9561, 281.9531, 281.9529, 281.958, 281.9629, 
    281.968, 281.9731, 281.978, 281.9832, 281.9883, 281.9932, 281.9983, 
    282.0034, 282.0083, 282.0134, 282.0186, 282.0356, 282.0527, 282.0696, 
    282.0867, 282.1035, 282.1206, 282.1375, 282.1545, 282.1714, 282.1885, 
    282.2056, 282.2224, 282.2395, 282.2559, 282.2722, 282.2883, 282.3044, 
    282.3208, 282.3369, 282.3533, 282.3694, 282.3857, 282.4019, 282.418, 
    282.4343, 282.4504, 282.4563, 282.4419, 282.4263, 282.4092, 282.3909, 
    282.3704, 282.3481, 282.3232, 282.2957, 282.2649, 282.2302, 282.1907, 
    282.1455, 282.094, 282.0911, 282.0879, 282.085, 282.082, 282.0789, 
    282.0759, 282.073, 282.0698, 282.0669, 282.064, 282.061, 282.0579, 
    282.0549, 282.0796, 282.1204, 282.165, 282.2146, 282.2698, 283.1794, 
    283.1895, 283.199, 283.208, 283.2168, 283.2251, 283.2329, 283.2405, 
    283.2505, 283.2659, 283.2812, 283.2966, 283.312, 283.3274, 283.3428, 
    283.3582, 283.3735, 283.3889, 283.4043, 283.4197, 283.4351, 283.4497, 
    283.4229, 283.396, 283.3691, 283.3425, 283.3157, 283.2888, 283.2622, 
    283.2354, 283.2085, 283.1816, 283.155, 283.1282, 283.1013, 283.0535, 
    282.9893, 282.916, 282.8313, 282.7324, 282.6157, 280.0166,
  281.7239, 281.9126, 282.1016, 282.2903, 282.479, 282.6677, 282.8567, 
    283.0454, 283.2341, 283.4229, 283.6116, 283.8005, 283.9453, 284.0068, 
    284.0681, 284.1294, 284.1907, 284.2522, 284.3135, 284.3748, 284.4363, 
    284.4976, 284.5588, 284.6201, 284.6816, 284.7415, 284.6819, 284.6221, 
    284.5623, 284.5027, 284.4429, 284.3831, 284.3235, 284.2637, 284.2039, 
    284.1443, 284.0845, 284.0247, 283.9651, 283.9431, 283.9392, 283.9353, 
    283.9314, 283.9275, 283.9236, 283.9197, 283.9158, 283.9119, 283.908, 
    283.9041, 283.9001, 283.8962, 283.9165, 283.9868, 284.0647, 284.1514, 
    284.248, 284.3567, 284.48, 284.6208, 287.4919, 287.6272, 287.7439, 
    287.8457, 287.9353, 288.0122, 287.8911, 287.77, 287.6489, 287.5278, 
    287.4067, 287.2856, 287.1646, 287.0435, 286.9224, 286.8013, 286.6802, 
    286.5591, 286.438, 286.3987, 286.3982, 286.3975, 286.397, 286.3965, 
    286.3958, 286.3953, 286.3948, 286.394, 286.3936, 286.3931, 286.3923, 
    286.3918, 286.4043, 286.4402, 286.4753, 286.5093, 286.5422, 286.5742, 
    286.6052, 286.6353, 286.6646, 286.6931, 286.7207, 286.7476, 286.7739, 
    286.7996, 286.8257, 286.8521, 286.8784, 286.9048, 286.9312, 286.9575, 
    286.9839, 287.01, 287.0364, 287.0627, 287.0891, 287.1155, 287.1418, 
    287.1138, 287.0601, 287.0066, 286.9529, 286.8992, 286.8457, 286.792, 
    286.7383, 286.6848, 286.6311, 286.5774, 286.5239, 286.4702, 286.4202, 
    286.3728, 286.3188, 286.2566, 286.1846, 286.0996, 285.998, 285.875, 
    285.7222, 285.5276, 285.2715, 284.9192, 283.637, 283.5906, 283.4612, 
    283.332, 283.2026, 283.0735, 282.9443, 282.8149, 282.6858, 282.5566, 
    282.4272, 282.2981, 282.1687, 282.0396, 281.9104, 281.8743, 281.8821, 
    281.8899, 281.8977, 281.9055, 281.9133, 281.9209, 281.9287, 281.9365, 
    281.9443, 281.9521, 281.96, 281.9678, 281.9739, 281.9771, 281.9805, 
    281.9836, 281.9868, 281.99, 281.9934, 281.9966, 281.9998, 282.0029, 
    282.0063, 282.0095, 282.0127, 282.0161, 282.0273, 282.0383, 282.0496, 
    282.0608, 282.072, 282.083, 282.0942, 282.1055, 282.1167, 282.1277, 
    282.1389, 282.1501, 282.1611, 282.1819, 282.2068, 282.2319, 282.2568, 
    282.2817, 282.3069, 282.3318, 282.3567, 282.3818, 282.4067, 282.4316, 
    282.4568, 282.4817, 282.4966, 282.4917, 282.4866, 282.4807, 282.4744, 
    282.467, 282.459, 283.0869, 283.114, 283.1372, 283.1572, 283.1746, 
    283.1899, 283.2034, 283.2024, 283.2014, 283.2007, 283.1997, 283.1987, 
    283.198, 283.197, 283.196, 283.1953, 283.1943, 283.1934, 283.1926, 
    283.1917, 283.1978, 283.2065, 283.2153, 283.2239, 283.2319, 283.24, 
    283.2478, 283.2554, 283.2627, 283.2698, 283.2766, 283.2834, 283.2898, 
    283.2988, 283.3123, 283.3257, 283.3391, 283.3525, 283.3662, 283.3796, 
    283.3931, 283.4065, 283.4199, 283.4336, 283.447, 283.4604, 283.4731, 
    283.4482, 283.4233, 283.3984, 283.3735, 283.3484, 283.3235, 283.2986, 
    283.2737, 283.2488, 283.2239, 283.1987, 283.1738, 283.1489, 283.1016, 
    283.0376, 282.9641, 282.8796, 282.781, 282.6643, 280.0681,
  281.9443, 282.135, 282.3254, 282.5161, 282.7068, 282.8975, 283.0879, 
    283.2786, 283.4692, 283.6599, 283.8503, 284.041, 284.1841, 284.2361, 
    284.2883, 284.3406, 284.3926, 284.4448, 284.4968, 284.5491, 284.6013, 
    284.6533, 284.7056, 284.7578, 284.8098, 284.8608, 284.7976, 284.7344, 
    284.6711, 284.6082, 284.5449, 284.4817, 284.4185, 284.3555, 284.2922, 
    284.229, 284.1658, 284.1025, 284.0396, 284.0134, 284.0051, 283.9968, 
    283.9885, 283.9802, 283.9719, 283.9636, 283.9553, 283.947, 283.9387, 
    283.9304, 283.9221, 283.9138, 283.9309, 284.002, 284.0818, 284.1726, 
    284.2769, 284.3972, 284.5381, 284.7056, 287.6614, 287.7866, 287.894, 
    287.9871, 288.0684, 288.1379, 288.0183, 287.8987, 287.7791, 287.6594, 
    287.54, 287.4204, 287.3008, 287.1812, 287.0615, 286.9419, 286.8223, 
    286.7026, 286.583, 286.5449, 286.5452, 286.5454, 286.5459, 286.5461, 
    286.5464, 286.5469, 286.5471, 286.5474, 286.5479, 286.5481, 286.5483, 
    286.5488, 286.562, 286.5994, 286.6362, 286.6729, 286.709, 286.7449, 
    286.7805, 286.8157, 286.8503, 286.885, 286.9192, 286.9531, 286.9866, 
    287.0195, 287.0291, 287.0386, 287.0479, 287.0574, 287.0669, 287.0762, 
    287.0857, 287.0952, 287.1047, 287.114, 287.1235, 287.1331, 287.1423, 
    287.1145, 287.0688, 287.0232, 286.9775, 286.9319, 286.8862, 286.8406, 
    286.7949, 286.7493, 286.7036, 286.658, 286.6123, 286.5667, 286.5217, 
    286.4741, 286.4199, 286.3574, 286.2849, 286.1995, 286.0977, 285.9739, 
    285.8203, 285.6248, 285.3672, 285.0132, 283.7244, 283.6775, 283.5325, 
    283.3875, 283.2427, 283.0977, 282.9526, 282.8076, 282.6626, 282.5176, 
    282.3728, 282.2278, 282.0828, 281.9377, 281.7927, 281.7593, 281.7778, 
    281.7964, 281.8149, 281.8335, 281.8521, 281.8708, 281.8894, 281.908, 
    281.9265, 281.9451, 281.9636, 281.9824, 281.9949, 281.9963, 281.9978, 
    281.9993, 282.0007, 282.002, 282.0034, 282.0049, 282.0063, 282.0078, 
    282.0093, 282.0105, 282.012, 282.0134, 282.0188, 282.0242, 282.0295, 
    282.0349, 282.0403, 282.0457, 282.051, 282.0564, 282.0618, 282.0669, 
    282.0723, 282.0776, 282.083, 282.1079, 282.1416, 282.1753, 282.209, 
    282.2429, 282.2766, 282.3103, 282.3442, 282.3779, 282.4116, 282.4456, 
    282.4792, 282.5129, 282.5369, 282.543, 282.5498, 282.5574, 282.5662, 
    282.5764, 282.5884, 283.155, 283.1807, 283.2021, 283.2207, 283.2366, 
    283.2507, 283.2627, 283.262, 283.2612, 283.2605, 283.2598, 283.2588, 
    283.2581, 283.2573, 283.2566, 283.2556, 283.2549, 283.2542, 283.2534, 
    283.2527, 283.2573, 283.2644, 283.2715, 283.2786, 283.2854, 283.2925, 
    283.2993, 283.3059, 283.3127, 283.3193, 283.3259, 283.3323, 283.3389, 
    283.3469, 283.3586, 283.3701, 283.3818, 283.3933, 283.4048, 283.4165, 
    283.428, 283.4397, 283.4512, 283.4626, 283.4744, 283.4858, 283.4968, 
    283.4739, 283.4507, 283.4275, 283.4045, 283.3813, 283.3582, 283.3352, 
    283.312, 283.2888, 283.2659, 283.2427, 283.2195, 283.1963, 283.1497, 
    283.0857, 283.0125, 282.928, 282.8293, 282.7129, 280.1199,
  282.0837, 282.2742, 282.4644, 282.6545, 282.8447, 283.0349, 283.2251, 
    283.4153, 283.6055, 283.7957, 283.9858, 284.176, 284.3154, 284.3582, 
    284.4009, 284.4436, 284.4866, 284.5293, 284.572, 284.6147, 284.6575, 
    284.7002, 284.7429, 284.7856, 284.8284, 284.8701, 284.8091, 284.748, 
    284.6873, 284.6262, 284.5654, 284.5044, 284.4436, 284.3826, 284.3215, 
    284.2607, 284.1997, 284.1389, 284.0779, 284.0518, 284.0422, 284.0325, 
    284.0227, 284.0129, 284.0029, 283.9929, 283.9829, 283.9729, 283.9626, 
    283.9521, 283.9419, 283.9314, 283.9478, 284.0215, 284.105, 284.2012, 
    284.3125, 284.4431, 284.5986, 284.7864, 287.5874, 287.7241, 287.8428, 
    287.9463, 288.0376, 288.1162, 288.0115, 287.9065, 287.8015, 287.6965, 
    287.5916, 287.4868, 287.3818, 287.2769, 287.1719, 287.0669, 286.9622, 
    286.8572, 286.7522, 286.7175, 286.7158, 286.7144, 286.7129, 286.7112, 
    286.7097, 286.7083, 286.7065, 286.7051, 286.7036, 286.7019, 286.7004, 
    286.699, 286.71, 286.7451, 286.7803, 286.8152, 286.8503, 286.8855, 
    286.9204, 286.9556, 286.9907, 287.0256, 287.0608, 287.0959, 287.1309, 
    287.1655, 287.1646, 287.1633, 287.1621, 287.1611, 287.1599, 287.1587, 
    287.1577, 287.1565, 287.1555, 287.1543, 287.1531, 287.1521, 287.1509, 
    287.1252, 287.0881, 287.0508, 287.0137, 286.9763, 286.9392, 286.9019, 
    286.8647, 286.8274, 286.7903, 286.7529, 286.7158, 286.6787, 286.6392, 
    286.592, 286.5383, 286.4766, 286.4048, 286.3201, 286.2192, 286.0967, 
    285.9446, 285.751, 285.4961, 285.1453, 283.8694, 283.8225, 283.6641, 
    283.5056, 283.3472, 283.1885, 283.03, 282.8716, 282.7131, 282.5544, 
    282.396, 282.2375, 282.0791, 281.9204, 281.762, 281.7261, 281.7473, 
    281.7688, 281.7903, 281.8118, 281.833, 281.8545, 281.876, 281.8972, 
    281.9187, 281.9402, 281.9614, 281.9829, 281.9968, 281.9968, 281.9971, 
    281.9971, 281.9971, 281.9971, 281.9971, 281.9971, 281.9971, 281.9971, 
    281.9971, 281.9971, 281.9971, 281.9973, 282.001, 282.0046, 282.0085, 
    282.0122, 282.0161, 282.0198, 282.0234, 282.0273, 282.031, 282.0347, 
    282.0386, 282.0422, 282.0459, 282.0725, 282.1099, 282.1475, 282.1853, 
    282.2236, 282.2622, 282.301, 282.3401, 282.3796, 282.4194, 282.4595, 
    282.5, 282.5408, 282.572, 282.5854, 282.6011, 282.6189, 282.6394, 
    282.6636, 282.6924, 283.249, 283.271, 283.2896, 283.3057, 283.3198, 
    283.3323, 283.343, 283.3403, 283.3376, 283.3347, 283.332, 283.3291, 
    283.3264, 283.3235, 283.3208, 283.3181, 283.3152, 283.3125, 283.3096, 
    283.3069, 283.3101, 283.3162, 283.3223, 283.3284, 283.3347, 283.3408, 
    283.3469, 283.353, 283.3591, 283.3652, 283.3713, 283.3774, 283.3835, 
    283.3914, 283.4019, 283.4126, 283.4233, 283.4341, 283.4448, 283.4556, 
    283.4661, 283.4768, 283.4875, 283.4983, 283.509, 283.5198, 283.5298, 
    283.5076, 283.4849, 283.4622, 283.4392, 283.4163, 283.3931, 283.3696, 
    283.3459, 283.322, 283.2981, 283.2739, 283.2495, 283.2249, 283.1758, 
    283.1089, 283.0327, 282.9448, 282.8428, 282.7222, 280.3049,
  282.1277, 282.3147, 282.5017, 282.689, 282.876, 283.0632, 283.2502, 
    283.4373, 283.6245, 283.8115, 283.9988, 284.1858, 284.3198, 284.353, 
    284.386, 284.4192, 284.4521, 284.4854, 284.5183, 284.5515, 284.5845, 
    284.6177, 284.6506, 284.6838, 284.7168, 284.749, 284.697, 284.645, 
    284.593, 284.5413, 284.4893, 284.4373, 284.3853, 284.3333, 284.2815, 
    284.2295, 284.1775, 284.1255, 284.0737, 284.0522, 284.0449, 284.0376, 
    284.03, 284.0222, 284.0144, 284.0061, 283.9978, 283.989, 283.9802, 
    283.9712, 283.9617, 283.9519, 283.9707, 284.0503, 284.1404, 284.2429, 
    284.3611, 284.4988, 284.6609, 284.855, 287.2832, 287.4475, 287.5935, 
    287.7241, 287.8418, 287.946, 287.8718, 287.7976, 287.7231, 287.6489, 
    287.5747, 287.5002, 287.426, 287.3518, 287.2773, 287.2031, 287.1289, 
    287.0544, 286.9802, 286.9519, 286.9456, 286.939, 286.9324, 286.9258, 
    286.9194, 286.9128, 286.9062, 286.8997, 286.8933, 286.8867, 286.8801, 
    286.8735, 286.8787, 286.905, 286.9316, 286.9583, 286.9849, 287.0115, 
    287.0381, 287.0645, 287.0911, 287.1177, 287.1443, 287.1709, 287.1975, 
    287.2236, 287.2195, 287.2151, 287.2109, 287.2068, 287.2024, 287.1982, 
    287.1938, 287.1897, 287.1855, 287.1812, 287.177, 287.1729, 287.1685, 
    287.1479, 287.1196, 287.0913, 287.0632, 287.0349, 287.0066, 286.9783, 
    286.95, 286.9219, 286.8936, 286.8652, 286.8369, 286.8086, 286.7756, 
    286.7297, 286.6775, 286.6174, 286.5474, 286.4653, 286.3672, 286.2478, 
    286.1001, 285.9119, 285.6638, 285.3228, 284.082, 284.0364, 283.8669, 
    283.6975, 283.5281, 283.3586, 283.1895, 283.02, 282.8506, 282.6812, 
    282.5117, 282.3423, 282.1729, 282.0034, 281.834, 281.79, 281.8049, 
    281.8196, 281.8342, 281.8491, 281.8638, 281.8787, 281.8933, 281.908, 
    281.9229, 281.9375, 281.9524, 281.967, 281.9763, 281.9753, 281.9746, 
    281.9736, 281.9727, 281.9719, 281.9709, 281.97, 281.9692, 281.9683, 
    281.9673, 281.9666, 281.9656, 281.9648, 281.9719, 281.979, 281.9863, 
    281.9934, 282.0005, 282.0076, 282.0149, 282.022, 282.0291, 282.0364, 
    282.0435, 282.0505, 282.0576, 282.0833, 282.1182, 282.1538, 282.1904, 
    282.228, 282.2666, 282.3064, 282.3472, 282.3892, 282.4321, 282.4766, 
    282.522, 282.5691, 282.606, 282.623, 282.6423, 282.6643, 282.6899, 
    282.7195, 282.7544, 283.3716, 283.3911, 283.4082, 283.4236, 283.4373, 
    283.4497, 283.4607, 283.4534, 283.446, 283.4387, 283.4314, 283.4241, 
    283.4167, 283.4097, 283.4023, 283.395, 283.3877, 283.3804, 283.373, 
    283.3657, 283.3667, 283.3716, 283.3762, 283.3811, 283.3857, 283.3906, 
    283.3953, 283.4001, 283.4048, 283.4097, 283.4143, 283.4192, 283.4238, 
    283.4309, 283.4419, 283.4529, 283.4639, 283.4751, 283.4861, 283.4971, 
    283.5081, 283.519, 283.53, 283.5413, 283.5522, 283.5632, 283.5737, 
    283.5515, 283.5286, 283.5051, 283.481, 283.4561, 283.4307, 283.4045, 
    283.3779, 283.3503, 283.3218, 283.2927, 283.2627, 283.2317, 283.1758, 
    283.1016, 283.0171, 282.9207, 282.8091, 282.6787, 280.6072,
  282.1714, 282.3555, 282.5393, 282.7234, 282.9075, 283.0916, 283.2754, 
    283.4595, 283.6436, 283.8276, 284.0115, 284.1956, 284.3245, 284.3479, 
    284.3711, 284.3945, 284.418, 284.4414, 284.4648, 284.4883, 284.5117, 
    284.5349, 284.5583, 284.5818, 284.6052, 284.6279, 284.585, 284.542, 
    284.499, 284.4561, 284.4131, 284.3701, 284.3271, 284.2842, 284.2412, 
    284.1982, 284.1553, 284.1123, 284.0693, 284.0525, 284.0479, 284.043, 
    284.0378, 284.0325, 284.0269, 284.021, 284.0149, 284.0083, 284.0015, 
    283.9944, 283.9868, 283.9788, 284.001, 284.0881, 284.186, 284.2969, 
    284.4233, 284.5691, 284.739, 284.9395, 287.0112, 287.1929, 287.3586, 
    287.5103, 287.6494, 287.7759, 287.7322, 287.6885, 287.6448, 287.6011, 
    287.5576, 287.5139, 287.4702, 287.4265, 287.3828, 287.3394, 287.2957, 
    287.252, 287.2083, 287.1865, 287.175, 287.1633, 287.1519, 287.1404, 
    287.1289, 287.1174, 287.106, 287.0945, 287.0828, 287.0713, 287.0598, 
    287.0483, 287.0471, 287.0652, 287.0833, 287.1013, 287.1194, 287.1375, 
    287.1555, 287.1736, 287.1917, 287.2097, 287.2278, 287.2458, 287.2639, 
    287.2817, 287.2744, 287.2668, 287.2595, 287.2522, 287.2449, 287.2375, 
    287.2302, 287.2229, 287.2156, 287.2083, 287.2009, 287.1936, 287.1863, 
    287.1707, 287.1514, 287.1321, 287.1128, 287.0935, 287.074, 287.0547, 
    287.0354, 287.0161, 286.9968, 286.9773, 286.958, 286.9387, 286.9119, 
    286.8672, 286.8167, 286.7581, 286.6902, 286.6104, 286.5149, 286.3992, 
    286.2556, 286.0725, 285.8318, 285.5005, 284.2947, 284.2502, 284.0698, 
    283.8896, 283.7092, 283.5291, 283.3486, 283.1685, 282.988, 282.8079, 
    282.6274, 282.447, 282.2668, 282.0864, 281.9062, 281.8542, 281.8623, 
    281.8704, 281.8784, 281.8865, 281.8945, 281.9026, 281.9106, 281.9187, 
    281.9268, 281.9348, 281.9431, 281.9512, 281.9558, 281.9539, 281.9521, 
    281.9502, 281.9485, 281.9465, 281.9448, 281.9431, 281.9412, 281.9395, 
    281.9375, 281.9358, 281.9338, 281.9324, 281.9429, 281.9534, 281.9639, 
    281.9746, 281.9851, 281.9956, 282.0061, 282.0166, 282.0273, 282.0378, 
    282.0483, 282.0588, 282.0693, 282.094, 282.1265, 282.1604, 282.1958, 
    282.2329, 282.2717, 282.3125, 282.3552, 282.4001, 282.4475, 282.4973, 
    282.55, 282.6057, 282.6504, 282.6719, 282.696, 282.7231, 282.7544, 
    282.7903, 282.832, 283.4775, 283.4985, 283.5173, 283.5347, 283.5505, 
    283.5652, 283.5781, 283.5662, 283.5544, 283.5427, 283.531, 283.519, 
    283.5073, 283.4956, 283.4836, 283.4719, 283.4602, 283.4482, 283.4365, 
    283.4248, 283.4233, 283.4268, 283.4302, 283.4336, 283.437, 283.4404, 
    283.4438, 283.4473, 283.4507, 283.4541, 283.4575, 283.4609, 283.4641, 
    283.4705, 283.4817, 283.4932, 283.5046, 283.5159, 283.5273, 283.5386, 
    283.55, 283.5613, 283.5728, 283.584, 283.5955, 283.6069, 283.6177, 
    283.5962, 283.5737, 283.55, 283.5256, 283.5, 283.4729, 283.4446, 283.415, 
    283.3838, 283.3508, 283.3162, 283.2795, 283.2407, 283.1758, 283.0918, 
    282.9971, 282.8894, 282.7661, 282.6238, 280.863,
  282.2151, 282.396, 282.5769, 282.7578, 282.9387, 283.1199, 283.3008, 
    283.4817, 283.6626, 283.8435, 284.0244, 284.2053, 284.3289, 284.3425, 
    284.3562, 284.3701, 284.3838, 284.3975, 284.4111, 284.425, 284.4387, 
    284.4524, 284.4661, 284.48, 284.4937, 284.5068, 284.4729, 284.439, 
    284.4048, 284.3708, 284.3369, 284.303, 284.269, 284.2349, 284.2009, 
    284.167, 284.1331, 284.0991, 284.0652, 284.0527, 284.0508, 284.0486, 
    284.0461, 284.0437, 284.0408, 284.0381, 284.0349, 284.0315, 284.0278, 
    284.0239, 284.0195, 284.0146, 284.0427, 284.1396, 284.2478, 284.3689, 
    284.5056, 284.6611, 284.8396, 285.0466, 286.7668, 286.9583, 287.137, 
    287.304, 287.4604, 287.6055, 287.5925, 287.5796, 287.5664, 287.5535, 
    287.5405, 287.5273, 287.5144, 287.5015, 287.4883, 287.4753, 287.4624, 
    287.4495, 287.4363, 287.4209, 287.4045, 287.3879, 287.3716, 287.355, 
    287.3386, 287.322, 287.3054, 287.2891, 287.2725, 287.2561, 287.2395, 
    287.2231, 287.2156, 287.2251, 287.2346, 287.2444, 287.2539, 287.2634, 
    287.2729, 287.2825, 287.292, 287.3018, 287.3113, 287.3208, 287.3303, 
    287.3396, 287.3293, 287.3188, 287.3083, 287.2979, 287.2874, 287.2771, 
    287.2666, 287.2561, 287.2456, 287.2354, 287.2249, 287.2144, 287.2039, 
    287.1936, 287.1831, 287.1726, 287.1624, 287.1519, 287.1416, 287.1311, 
    287.1206, 287.1104, 287.0999, 287.0896, 287.0791, 287.0688, 287.0481, 
    287.0049, 286.9556, 286.8989, 286.833, 286.7554, 286.6628, 286.5505, 
    286.4109, 286.2334, 285.9995, 285.678, 284.5076, 284.4641, 284.2727, 
    284.0815, 283.8904, 283.6992, 283.5081, 283.3169, 283.1255, 282.9343, 
    282.7432, 282.552, 282.3608, 282.1694, 281.9783, 281.9182, 281.9197, 
    281.9211, 281.9226, 281.9238, 281.9253, 281.9268, 281.9282, 281.9294, 
    281.9309, 281.9324, 281.9338, 281.9351, 281.9351, 281.9324, 281.9297, 
    281.927, 281.9241, 281.9214, 281.9187, 281.916, 281.9133, 281.9106, 
    281.9077, 281.905, 281.9023, 281.8999, 281.9138, 281.9277, 281.9417, 
    281.9556, 281.9695, 281.9834, 281.9976, 282.0115, 282.0254, 282.0393, 
    282.0532, 282.0671, 282.0811, 282.105, 282.1353, 282.1672, 282.2017, 
    282.238, 282.2773, 282.3193, 282.3645, 282.4133, 282.4663, 282.5237, 
    282.5862, 282.6548, 282.7117, 282.7385, 282.7683, 282.802, 282.8396, 
    282.8826, 282.9319, 283.5703, 283.5952, 283.6182, 283.6396, 283.6597, 
    283.6785, 283.6956, 283.6792, 283.6628, 283.6467, 283.6304, 283.614, 
    283.5977, 283.5815, 283.5652, 283.5488, 283.5325, 283.5164, 283.5, 
    283.4836, 283.48, 283.4819, 283.4841, 283.4861, 283.488, 283.4902, 
    283.4922, 283.4944, 283.4963, 283.4983, 283.5005, 283.5024, 283.5046, 
    283.51, 283.5217, 283.5334, 283.5452, 283.5569, 283.5686, 283.5803, 
    283.5918, 283.6035, 283.6152, 283.627, 283.6387, 283.6504, 283.6616, 
    283.6416, 283.6204, 283.5979, 283.5737, 283.5481, 283.5205, 283.4907, 
    283.4587, 283.4243, 283.387, 283.3462, 283.3018, 283.2532, 283.1758, 
    283.0784, 282.9697, 282.8477, 282.7097, 282.552, 281.0825,
  282.2588, 282.4368, 282.6145, 282.7925, 282.9702, 283.1482, 283.3259, 
    283.5039, 283.6816, 283.8596, 284.0374, 284.2153, 284.3333, 284.3374, 
    284.3413, 284.3455, 284.3496, 284.3535, 284.3577, 284.3618, 284.3657, 
    284.3699, 284.374, 284.3779, 284.3821, 284.3857, 284.3608, 284.3357, 
    284.3108, 284.2859, 284.2607, 284.2358, 284.2107, 284.1858, 284.1609, 
    284.1357, 284.1108, 284.0857, 284.0608, 284.0532, 284.0537, 284.0544, 
    284.0549, 284.0557, 284.0566, 284.0576, 284.0586, 284.0596, 284.061, 
    284.0623, 284.064, 284.0659, 284.103, 284.2139, 284.3357, 284.4702, 
    284.6199, 284.7866, 284.9744, 285.1868, 286.5457, 286.741, 286.9272, 
    287.105, 287.2747, 287.4353, 287.4529, 287.4705, 287.4883, 287.5059, 
    287.5234, 287.541, 287.5586, 287.5762, 287.594, 287.6116, 287.6292, 
    287.6467, 287.6643, 287.6555, 287.634, 287.6125, 287.5911, 287.5696, 
    287.5481, 287.5266, 287.5051, 287.4836, 287.4622, 287.4407, 287.4192, 
    287.3977, 287.384, 287.3853, 287.3862, 287.3872, 287.3884, 287.3894, 
    287.3904, 287.3916, 287.3926, 287.3936, 287.3948, 287.3958, 287.3967, 
    287.3977, 287.3843, 287.3706, 287.3572, 287.3435, 287.3301, 287.3164, 
    287.303, 287.2893, 287.2759, 287.2622, 287.2488, 287.2351, 287.2217, 
    287.2163, 287.2148, 287.2134, 287.2119, 287.2104, 287.209, 287.2075, 
    287.2061, 287.2046, 287.2031, 287.2017, 287.2002, 287.1987, 287.1846, 
    287.1426, 287.0947, 287.0398, 286.9758, 286.9006, 286.8108, 286.7017, 
    286.5664, 286.3943, 286.1675, 285.8555, 284.7202, 284.6777, 284.4758, 
    284.2737, 284.0715, 283.8694, 283.6672, 283.4651, 283.2632, 283.061, 
    282.8589, 282.6567, 282.4546, 282.2524, 282.0505, 281.9824, 281.9771, 
    281.9719, 281.9666, 281.9614, 281.9561, 281.9507, 281.9456, 281.9402, 
    281.9351, 281.9297, 281.9246, 281.9192, 281.9146, 281.9109, 281.9072, 
    281.9036, 281.8999, 281.8962, 281.8926, 281.8889, 281.8853, 281.8816, 
    281.8779, 281.8743, 281.8706, 281.8674, 281.8848, 281.9021, 281.9194, 
    281.9368, 281.9541, 281.9714, 281.9888, 282.0061, 282.0234, 282.0408, 
    282.0581, 282.0754, 282.0928, 282.1162, 282.1443, 282.1746, 282.2078, 
    282.2439, 282.2834, 282.3274, 282.3757, 282.4297, 282.49, 282.5581, 
    282.6357, 282.7246, 282.801, 282.8347, 282.8716, 282.9126, 282.958, 
    283.0088, 283.0657, 283.6523, 283.6826, 283.7114, 283.7388, 283.7649, 
    283.7898, 283.813, 283.7922, 283.7715, 283.7507, 283.7297, 283.709, 
    283.6882, 283.6675, 283.6467, 283.6257, 283.605, 283.5842, 283.5635, 
    283.5427, 283.5366, 283.5371, 283.5378, 283.5386, 283.5393, 283.54, 
    283.5408, 283.5415, 283.5422, 283.5427, 283.5435, 283.5442, 283.5449, 
    283.5496, 283.5615, 283.5737, 283.5857, 283.5977, 283.6099, 283.6218, 
    283.6338, 283.6458, 283.658, 283.6699, 283.6819, 283.6941, 283.7056, 
    283.688, 283.6689, 283.6484, 283.6257, 283.6013, 283.5742, 283.5444, 
    283.5112, 283.4744, 283.4329, 283.386, 283.3323, 283.2708, 283.1758, 
    283.0593, 282.9312, 282.7896, 282.6316, 282.4551, 281.2729,
  282.3025, 282.4773, 282.6521, 282.8269, 283.0017, 283.1765, 283.3511, 
    283.5259, 283.7007, 283.8755, 284.0503, 284.2251, 284.3376, 284.332, 
    284.3264, 284.3208, 284.3154, 284.3098, 284.3042, 284.2986, 284.293, 
    284.2874, 284.2817, 284.2761, 284.2705, 284.2646, 284.2488, 284.2327, 
    284.2166, 284.2007, 284.1846, 284.1687, 284.1526, 284.1365, 284.1206, 
    284.1045, 284.0886, 284.0725, 284.0564, 284.0535, 284.0569, 284.0605, 
    284.0647, 284.0693, 284.0745, 284.0803, 284.0872, 284.095, 284.104, 
    284.1147, 284.1279, 284.144, 284.1995, 284.3303, 284.4712, 284.6235, 
    284.7886, 284.9678, 285.1636, 285.3782, 286.3445, 286.5393, 286.7288, 
    286.9131, 287.0923, 287.2651, 287.3132, 287.3616, 287.4099, 287.458, 
    287.5063, 287.5547, 287.6028, 287.6511, 287.6995, 287.7476, 287.7959, 
    287.8442, 287.8923, 287.8899, 287.8635, 287.8369, 287.8105, 287.7842, 
    287.7576, 287.7312, 287.7048, 287.6782, 287.6519, 287.6255, 287.5989, 
    287.5725, 287.5527, 287.5452, 287.5378, 287.5303, 287.5229, 287.5154, 
    287.5081, 287.5005, 287.4932, 287.4856, 287.4783, 287.4707, 287.4634, 
    287.4558, 287.4392, 287.4224, 287.4058, 287.3892, 287.3726, 287.3557, 
    287.3391, 287.3225, 287.3059, 287.2893, 287.2725, 287.2559, 287.2393, 
    287.239, 287.2466, 287.2539, 287.2615, 287.269, 287.2764, 287.2839, 
    287.2915, 287.2988, 287.3064, 287.314, 287.3213, 287.3289, 287.3208, 
    287.28, 287.2339, 287.1804, 287.1187, 287.0457, 286.9587, 286.853, 
    286.7219, 286.5549, 286.3352, 286.033, 284.9331, 284.8916, 284.6787, 
    284.4656, 284.2527, 284.0396, 283.8267, 283.6135, 283.4006, 283.1875, 
    282.9746, 282.7615, 282.5486, 282.3357, 282.1226, 282.0464, 282.0347, 
    282.0227, 282.0107, 281.9988, 281.9868, 281.9749, 281.9629, 281.9509, 
    281.939, 281.9272, 281.9153, 281.9033, 281.8938, 281.8894, 281.8848, 
    281.8801, 281.8757, 281.8711, 281.8665, 281.8621, 281.8574, 281.8528, 
    281.8481, 281.8438, 281.8391, 281.835, 281.8557, 281.8765, 281.8972, 
    281.918, 281.9387, 281.9595, 281.98, 282.0007, 282.0215, 282.0422, 
    282.063, 282.0837, 282.1045, 282.1274, 282.1536, 282.1824, 282.2144, 
    282.2502, 282.2908, 282.3367, 282.3892, 282.45, 282.521, 282.6052, 
    282.7068, 282.8313, 282.9429, 282.9851, 283.0305, 283.0796, 283.1328, 
    283.1907, 283.2539, 283.7251, 283.762, 283.7979, 283.8325, 283.8665, 
    283.8994, 283.9304, 283.9053, 283.8799, 283.8545, 283.8293, 283.804, 
    283.7788, 283.7534, 283.728, 283.7029, 283.6775, 283.6521, 283.627, 
    283.6016, 283.593, 283.5925, 283.5918, 283.5911, 283.5906, 283.5898, 
    283.5891, 283.5886, 283.5879, 283.5872, 283.5867, 283.5859, 283.5852, 
    283.5891, 283.6016, 283.6138, 283.6262, 283.6387, 283.6509, 283.6633, 
    283.6758, 283.688, 283.7004, 283.7129, 283.7251, 283.7375, 283.7495, 
    283.7351, 283.7192, 283.7019, 283.6824, 283.6604, 283.6357, 283.6074, 
    283.5752, 283.5376, 283.4934, 283.4409, 283.3772, 283.2986, 283.1758, 
    283.0298, 282.8723, 282.7021, 282.5173, 282.3162, 281.4395,
  282.3462, 282.5181, 282.6897, 282.8613, 283.033, 283.2046, 283.3765, 
    283.5481, 283.7197, 283.8914, 284.0632, 284.2349, 284.3423, 284.3269, 
    284.3115, 284.2964, 284.281, 284.2659, 284.2505, 284.2354, 284.22, 
    284.2046, 284.1895, 284.1741, 284.1589, 284.1436, 284.1367, 284.1296, 
    284.1226, 284.1155, 284.1084, 284.1016, 284.0945, 284.0874, 284.0803, 
    284.0732, 284.0664, 284.0593, 284.0522, 284.0537, 284.0601, 284.0669, 
    284.075, 284.0842, 284.0947, 284.1072, 284.1221, 284.1401, 284.1624, 
    284.1907, 284.2275, 284.2781, 284.3772, 284.5391, 284.707, 284.8818, 
    285.0635, 285.2524, 285.4495, 285.6548, 286.1611, 286.3518, 286.5405, 
    286.7275, 286.9126, 287.0947, 287.1736, 287.2527, 287.3315, 287.4104, 
    287.4893, 287.5681, 287.647, 287.7261, 287.8049, 287.8838, 287.9626, 
    288.0415, 288.1204, 288.1245, 288.093, 288.0615, 288.03, 287.9988, 
    287.9673, 287.9358, 287.9043, 287.873, 287.8416, 287.8101, 287.7786, 
    287.7473, 287.7212, 287.7051, 287.6892, 287.6733, 287.6575, 287.6414, 
    287.6255, 287.6096, 287.5935, 287.5776, 287.5618, 287.5457, 287.5298, 
    287.5137, 287.4941, 287.4744, 287.4546, 287.4348, 287.415, 287.3953, 
    287.3755, 287.3557, 287.3359, 287.3162, 287.2964, 287.2766, 287.2568, 
    287.2617, 287.2781, 287.2947, 287.311, 287.3274, 287.344, 287.3604, 
    287.3767, 287.3931, 287.4097, 287.426, 287.4424, 287.459, 287.457, 
    287.4177, 287.3728, 287.3213, 287.2612, 287.1909, 287.1067, 287.0044, 
    286.8774, 286.7158, 286.5032, 286.2104, 285.1458, 285.1055, 284.8816, 
    284.6577, 284.4338, 284.21, 283.9858, 283.762, 283.5381, 283.3142, 
    283.0903, 282.8665, 282.6426, 282.4187, 282.1946, 282.1106, 282.092, 
    282.0735, 282.0547, 282.0361, 282.0176, 281.999, 281.9805, 281.9617, 
    281.9431, 281.9246, 281.906, 281.8875, 281.8733, 281.8679, 281.8623, 
    281.8569, 281.8513, 281.8459, 281.8403, 281.835, 281.8293, 281.824, 
    281.8184, 281.813, 281.8076, 281.8025, 281.8267, 281.8508, 281.8748, 
    281.8989, 281.9231, 281.9473, 281.9714, 281.9956, 282.0198, 282.0437, 
    282.0679, 282.092, 282.1162, 282.1389, 282.1631, 282.1904, 282.2214, 
    282.2573, 282.2988, 282.3474, 282.4055, 282.4758, 282.5627, 282.6731, 
    282.8176, 283.0149, 283.2046, 283.2549, 283.3071, 283.3613, 283.418, 
    283.4766, 283.5378, 283.7903, 283.8345, 283.8784, 283.9216, 283.9646, 
    284.0071, 284.0481, 284.0181, 283.9883, 283.9585, 283.9287, 283.8989, 
    283.8691, 283.8394, 283.8096, 283.7798, 283.75, 283.7202, 283.6904, 
    283.6606, 283.6497, 283.6477, 283.6458, 283.6438, 283.6416, 283.6396, 
    283.6377, 283.6357, 283.6335, 283.6316, 283.6296, 283.6277, 283.6255, 
    283.6287, 283.6414, 283.6541, 283.6667, 283.6794, 283.6921, 283.7048, 
    283.7175, 283.7302, 283.7429, 283.7559, 283.7686, 283.7812, 283.7935, 
    283.7832, 283.7717, 283.7585, 283.7437, 283.7266, 283.7065, 283.6831, 
    283.6548, 283.6204, 283.5774, 283.5225, 283.4495, 283.3481, 283.1755, 
    282.9771, 282.7708, 282.5564, 282.3333, 282.1011, 281.5864,
  282.4463, 282.6086, 282.7712, 282.9336, 283.0959, 283.2583, 283.4207, 
    283.5833, 283.7456, 283.908, 284.0703, 284.2305, 284.3289, 284.3098, 
    284.2908, 284.2717, 284.2527, 284.2334, 284.2144, 284.1953, 284.1763, 
    284.1572, 284.1382, 284.1228, 284.1108, 284.0991, 284.105, 284.1108, 
    284.1167, 284.1226, 284.1284, 284.134, 284.1399, 284.1458, 284.1516, 
    284.1575, 284.1497, 284.1418, 284.1338, 284.1348, 284.1404, 284.147, 
    284.1545, 284.1636, 284.5273, 284.5439, 284.5576, 284.5688, 284.5813, 
    284.5942, 284.6055, 284.6157, 284.6853, 284.8701, 285.0549, 285.2397, 
    285.4243, 285.6091, 285.7939, 285.9788, 286.1636, 286.3408, 286.5183, 
    286.6956, 286.873, 287.0493, 287.1416, 287.2339, 287.3262, 287.4185, 
    287.5107, 287.6028, 287.6951, 287.7861, 287.8755, 287.9651, 288.0547, 
    288.144, 288.2336, 288.2397, 288.2065, 288.1733, 288.1404, 288.1072, 
    288.074, 288.0408, 288.0085, 287.9761, 287.9438, 287.9114, 287.8792, 
    287.8469, 287.8188, 287.7993, 287.7795, 287.76, 287.7402, 287.7205, 
    287.7007, 287.6807, 287.6606, 287.6406, 287.6206, 287.6006, 287.5806, 
    287.5605, 287.5398, 287.519, 287.4983, 287.4775, 287.457, 287.436, 
    287.4153, 287.3945, 287.3738, 287.3528, 287.332, 287.3113, 287.2905, 
    287.2971, 287.3167, 287.3364, 287.356, 287.3748, 287.3928, 287.4106, 
    287.4287, 287.4468, 287.4646, 287.4827, 287.5005, 287.5186, 287.5176, 
    287.478, 287.4333, 287.3826, 287.3232, 287.2537, 287.1709, 287.0703, 
    286.9463, 286.7891, 286.583, 286.3018, 285.1924, 285.1487, 284.9216, 
    284.696, 284.4709, 284.2451, 284.0193, 283.7935, 283.5676, 283.3416, 
    283.1157, 282.8899, 282.6641, 282.438, 282.2122, 282.1191, 282.0884, 
    282.0706, 282.0527, 282.0352, 282.0173, 281.9998, 281.9819, 281.9641, 
    281.9465, 281.9287, 281.9109, 281.8933, 281.8809, 281.8772, 281.8721, 
    281.8669, 281.8618, 281.8569, 281.8518, 281.8467, 281.8416, 281.8364, 
    281.8315, 281.8264, 281.8213, 281.8167, 281.8391, 281.8613, 281.8838, 
    281.9062, 281.9285, 281.9509, 281.9731, 281.9956, 282.0181, 282.0403, 
    282.0627, 282.085, 282.1089, 282.1304, 282.1526, 282.1777, 282.2068, 
    282.2407, 282.281, 282.3293, 282.3887, 282.4631, 282.5591, 282.688, 
    283.3242, 283.3628, 283.4053, 283.4612, 283.5171, 283.5732, 283.6292, 
    283.6851, 283.7412, 283.7971, 283.853, 283.9092, 283.9651, 284.0161, 
    284.062, 284.1067, 284.0764, 284.0464, 284.0161, 283.9861, 283.9558, 
    283.9258, 283.8955, 283.8652, 283.8352, 283.8049, 283.7754, 283.7458, 
    283.7161, 283.7053, 283.7036, 283.7017, 283.7, 283.698, 283.696, 
    283.6943, 283.6924, 283.6904, 283.6873, 283.6826, 283.678, 283.6733, 
    283.6741, 283.6841, 283.6941, 283.7043, 283.7144, 283.7244, 283.7346, 
    283.7446, 283.7546, 283.7646, 283.7749, 283.7852, 283.7954, 283.8054, 
    283.7952, 283.7837, 283.7705, 283.3201, 283.2937, 283.2727, 283.2556, 
    283.2427, 283.2329, 283.2246, 283.2173, 283.2109, 283.2051, 283.0371, 
    282.7937, 282.5503, 282.3069, 282.0635, 281.8201, 281.5767,
  282.6213, 282.7664, 282.9111, 283.0559, 283.2009, 283.3457, 283.4907, 
    283.6355, 283.7803, 283.9253, 284.0701, 284.207, 284.2917, 284.2766, 
    284.2617, 284.2466, 284.2317, 284.2166, 284.2017, 284.1865, 284.1716, 
    284.1565, 284.1416, 284.1384, 284.1472, 284.1562, 284.1802, 284.2041, 
    284.228, 284.252, 284.2759, 284.2998, 284.3237, 284.3474, 284.3713, 
    284.3953, 284.3765, 284.3574, 284.3376, 284.332, 284.3333, 284.3347, 
    284.3367, 284.3386, 284.7874, 284.7964, 284.8037, 284.8098, 284.8254, 
    284.8486, 284.8696, 284.8884, 284.9617, 285.1411, 285.3203, 285.4998, 
    285.6792, 285.8586, 286.0381, 286.2173, 286.3967, 286.5518, 286.7065, 
    286.8613, 287.0161, 287.1702, 287.2527, 287.3354, 287.418, 287.5005, 
    287.5833, 287.6658, 287.7483, 287.8264, 287.8999, 287.9734, 288.0469, 
    288.1204, 288.1938, 288.1968, 288.166, 288.1355, 288.1047, 288.0742, 
    288.0437, 288.0129, 287.9854, 287.9575, 287.9297, 287.9021, 287.8743, 
    287.8464, 287.8225, 287.8054, 287.7883, 287.7715, 287.7544, 287.7373, 
    287.7197, 287.7014, 287.6833, 287.665, 287.647, 287.6287, 287.6104, 
    287.5923, 287.5735, 287.5544, 287.5356, 287.5168, 287.498, 287.479, 
    287.46, 287.4407, 287.4216, 287.4026, 287.3833, 287.3643, 287.3452, 
    287.3494, 287.3645, 287.3796, 287.395, 287.4072, 287.417, 287.4268, 
    287.4363, 287.446, 287.4556, 287.4653, 287.4749, 287.4846, 287.4775, 
    287.4363, 287.3909, 287.3401, 287.2798, 287.2097, 287.1265, 287.0261, 
    286.9031, 286.7485, 286.5488, 286.2803, 285.011, 284.959, 284.741, 
    284.5288, 284.3169, 284.1008, 283.8848, 283.6689, 283.4529, 283.2371, 
    283.021, 282.8049, 282.5891, 282.373, 282.1572, 282.054, 282.0034, 
    281.9966, 281.9897, 281.9829, 281.9761, 281.9692, 281.9624, 281.9556, 
    281.9487, 281.9419, 281.9351, 281.9282, 281.926, 281.9275, 281.9248, 
    281.9219, 281.9189, 281.916, 281.9131, 281.9102, 281.9072, 281.9043, 
    281.9014, 281.8984, 281.8955, 281.8931, 281.9067, 281.9204, 281.9343, 
    281.948, 281.9617, 281.9753, 281.989, 282.0029, 282.0166, 282.0303, 
    282.0439, 282.0576, 282.0762, 282.0952, 282.1143, 282.136, 282.1611, 
    282.1907, 282.2261, 282.2686, 282.321, 282.3872, 282.4736, 282.5911, 
    283.0825, 283.1533, 283.2214, 283.2944, 283.3677, 283.4407, 283.5139, 
    283.5869, 283.6602, 283.7332, 283.8064, 283.8794, 283.9526, 284.009, 
    284.0483, 284.0869, 284.062, 284.0369, 284.012, 283.9871, 283.9619, 
    283.937, 283.9119, 283.887, 283.8621, 283.8369, 283.8137, 283.7905, 
    283.7671, 283.76, 283.7603, 283.7605, 283.7607, 283.7612, 283.7615, 
    283.7617, 283.762, 283.7622, 283.7581, 283.749, 283.7402, 283.7312, 
    283.7266, 283.7302, 283.7339, 283.7373, 283.741, 283.7446, 283.748, 
    283.7517, 283.7551, 283.7585, 283.762, 283.7654, 283.769, 283.7725, 
    283.7556, 283.7363, 283.7141, 282.9626, 282.9421, 282.9255, 282.9119, 
    282.9014, 282.8933, 282.886, 282.8794, 282.8735, 282.8682, 282.7141, 
    282.491, 282.2678, 282.0447, 281.8215, 281.5984, 281.3752,
  282.7964, 282.9238, 283.051, 283.1785, 283.3059, 283.4331, 283.5605, 
    283.6877, 283.8152, 283.9426, 284.0698, 284.1838, 284.2546, 284.2437, 
    284.2327, 284.2217, 284.2107, 284.1997, 284.1887, 284.178, 284.167, 
    284.156, 284.145, 284.1543, 284.1838, 284.2136, 284.2556, 284.2976, 
    284.3394, 284.3813, 284.4233, 284.4653, 284.5073, 284.5493, 284.5911, 
    284.6331, 284.6077, 284.5811, 284.5532, 284.5427, 284.5408, 284.5381, 
    284.5354, 284.5317, 285.0193, 285.0234, 285.0269, 285.0298, 285.0518, 
    285.0903, 285.1255, 285.158, 285.2378, 285.4119, 285.5859, 285.76, 
    285.9341, 286.1082, 286.282, 286.4561, 286.6301, 286.7625, 286.8948, 
    287.0271, 287.1594, 287.291, 287.364, 287.4368, 287.5098, 287.5828, 
    287.6558, 287.7288, 287.8018, 287.8669, 287.9243, 287.9817, 288.0393, 
    288.0967, 288.1543, 288.1536, 288.1255, 288.0974, 288.0693, 288.0415, 
    288.0134, 287.9854, 287.9622, 287.939, 287.9158, 287.8926, 287.8694, 
    287.8462, 287.8259, 287.8118, 287.7974, 287.783, 287.7686, 287.7542, 
    287.7388, 287.7224, 287.7061, 287.6895, 287.6731, 287.6567, 287.6404, 
    287.6238, 287.6069, 287.5901, 287.5732, 287.5562, 287.5393, 287.522, 
    287.5044, 287.4871, 287.4695, 287.4521, 287.4348, 287.4172, 287.3999, 
    287.4016, 287.4124, 287.4231, 287.4338, 287.4399, 287.4412, 287.4426, 
    287.4438, 287.4453, 287.4465, 287.448, 287.4492, 287.4507, 287.4377, 
    287.3958, 287.3501, 287.3003, 287.2395, 287.1689, 287.0854, 286.9856, 
    286.864, 286.7124, 286.5186, 286.2615, 284.8203, 284.76, 284.5554, 
    284.3601, 284.1626, 283.9565, 283.7505, 283.5444, 283.3384, 283.1323, 
    282.9263, 282.7202, 282.5142, 282.3081, 282.1021, 281.9885, 281.9185, 
    281.9226, 281.9265, 281.9307, 281.9348, 281.9387, 281.9429, 281.947, 
    281.9509, 281.9551, 281.9592, 281.9631, 281.9709, 281.978, 281.9773, 
    281.9766, 281.9758, 281.9751, 281.9744, 281.9736, 281.9729, 281.9722, 
    281.9714, 281.9707, 281.9697, 281.9695, 281.9746, 281.9795, 281.9846, 
    281.9897, 281.9949, 281.9998, 282.0049, 282.01, 282.0151, 282.0203, 
    282.0251, 282.0303, 282.043, 282.0593, 282.0752, 282.0933, 282.1145, 
    282.1394, 282.1692, 282.2053, 282.2502, 282.3071, 282.3823, 282.4858, 
    282.8479, 282.946, 283.0376, 283.1279, 283.218, 283.3083, 283.3987, 
    283.4888, 283.5791, 283.6694, 283.7595, 283.8499, 283.9402, 284.0017, 
    284.0349, 284.0674, 284.0474, 284.0276, 284.0078, 283.988, 283.968, 
    283.9482, 283.9285, 283.9087, 283.8887, 283.8689, 283.8521, 283.8352, 
    283.8181, 283.8145, 283.8169, 283.8193, 283.8218, 283.8242, 283.8267, 
    283.8291, 283.8315, 283.834, 283.8286, 283.8154, 283.8022, 283.7891, 
    283.7793, 283.7764, 283.7734, 283.7705, 283.7676, 283.7646, 283.7617, 
    283.7588, 283.7556, 283.7522, 283.7485, 283.7446, 283.7405, 283.7361, 
    283.7117, 283.6833, 283.6501, 282.6663, 282.6453, 282.6284, 282.614, 
    282.5994, 282.5835, 282.5693, 282.5562, 282.5442, 282.5332, 282.3911, 
    282.1882, 281.9854, 281.7825, 281.5798, 281.377, 281.1741,
  282.9714, 283.0813, 283.1912, 283.3008, 283.4106, 283.5205, 283.6304, 
    283.7402, 283.8501, 283.9597, 284.0696, 284.1604, 284.2175, 284.2107, 
    284.2036, 284.1968, 284.1899, 284.1829, 284.176, 284.1692, 284.1621, 
    284.1553, 284.1484, 284.1702, 284.2205, 284.2708, 284.3308, 284.3909, 
    284.4509, 284.511, 284.5708, 284.6309, 284.6909, 284.751, 284.8108, 
    284.8708, 284.8433, 284.8137, 284.782, 284.7688, 284.7644, 284.7593, 
    284.7532, 284.7458, 285.2275, 285.229, 285.2302, 285.2312, 285.2622, 
    285.3198, 285.3738, 285.4246, 285.5142, 285.6829, 285.8516, 286.02, 
    286.1887, 286.3574, 286.5261, 286.6948, 286.8635, 286.9731, 287.083, 
    287.1929, 287.3025, 287.4116, 287.4751, 287.5383, 287.6016, 287.665, 
    287.7283, 287.7915, 287.855, 287.9072, 287.9487, 287.9902, 288.0315, 
    288.073, 288.1145, 288.1104, 288.085, 288.0596, 288.0339, 288.0085, 
    287.9832, 287.9575, 287.939, 287.9204, 287.9016, 287.8831, 287.8645, 
    287.8459, 287.8296, 287.8179, 287.8062, 287.7944, 287.7827, 287.771, 
    287.7578, 287.7432, 287.7285, 287.7139, 287.6995, 287.6848, 287.6702, 
    287.6555, 287.6406, 287.6255, 287.6106, 287.5955, 287.5806, 287.5647, 
    287.5491, 287.5332, 287.5176, 287.5017, 287.4861, 287.4702, 287.4546, 
    287.4539, 287.46, 287.4663, 287.4727, 287.4724, 287.4653, 287.4585, 
    287.4514, 287.4446, 287.4375, 287.4307, 287.4236, 287.4167, 287.3982, 
    287.356, 287.311, 287.2632, 287.2019, 287.1309, 287.0476, 286.9482, 
    286.8281, 286.6797, 286.4912, 286.2449, 284.6191, 284.551, 284.3645, 
    284.1897, 284.0083, 283.8123, 283.6162, 283.4199, 283.2239, 283.0276, 
    282.8315, 282.6353, 282.4392, 282.2432, 282.0469, 281.9233, 281.8335, 
    281.8484, 281.8635, 281.8784, 281.8933, 281.9084, 281.9233, 281.9382, 
    281.9534, 281.9683, 281.9832, 281.9983, 282.0161, 282.0286, 282.0298, 
    282.0312, 282.0327, 282.0342, 282.0356, 282.0371, 282.0383, 282.0398, 
    282.0413, 282.0427, 282.0442, 282.0459, 282.0422, 282.0386, 282.0352, 
    282.0315, 282.0278, 282.0244, 282.0208, 282.0173, 282.0137, 282.01, 
    282.0066, 282.0029, 282.0095, 282.0227, 282.0354, 282.0498, 282.0667, 
    282.0864, 282.1104, 282.1396, 282.176, 282.2227, 282.2849, 282.3716, 
    282.6201, 282.7415, 282.8538, 282.9612, 283.0686, 283.1758, 283.2832, 
    283.3906, 283.498, 283.6055, 283.7129, 283.8203, 283.9275, 283.9946, 
    284.0215, 284.0476, 284.033, 284.0183, 284.0037, 283.989, 283.9744, 
    283.9597, 283.9448, 283.9302, 283.9155, 283.9009, 283.8904, 283.8799, 
    283.8691, 283.8691, 283.8735, 283.8782, 283.8828, 283.8875, 283.8921, 
    283.8967, 283.9011, 283.9058, 283.8994, 283.8818, 283.8643, 283.8469, 
    283.832, 283.8228, 283.8132, 283.8037, 283.7942, 283.7847, 283.7751, 
    283.7656, 283.7563, 283.7458, 283.7346, 283.7227, 283.7097, 283.6958, 
    283.6624, 283.6233, 283.5769, 282.4167, 282.3916, 282.3708, 282.3535, 
    282.3298, 282.3003, 282.2725, 282.2468, 282.2224, 282.2, 282.0681, 
    281.8855, 281.7029, 281.5205, 281.3379, 281.1553, 280.9729,
  283.1465, 283.2388, 283.3311, 283.4233, 283.5156, 283.6079, 283.7002, 
    283.7925, 283.8848, 283.9771, 284.0693, 284.137, 284.1804, 284.1775, 
    284.1748, 284.1719, 284.1689, 284.166, 284.1633, 284.1604, 284.1575, 
    284.1545, 284.1519, 284.1858, 284.2568, 284.3281, 284.4062, 284.4841, 
    284.5623, 284.6404, 284.7185, 284.7964, 284.8745, 284.9526, 285.0308, 
    285.1086, 285.0833, 285.0554, 285.0249, 285.0115, 285.0066, 285.0005, 
    284.9934, 284.9846, 285.4155, 285.416, 285.4163, 285.4167, 285.4583, 
    285.5386, 285.615, 285.688, 285.7903, 285.9536, 286.1169, 286.2803, 
    286.4436, 286.6069, 286.7703, 286.9336, 287.0969, 287.1841, 287.2712, 
    287.3584, 287.4458, 287.5325, 287.5862, 287.6399, 287.6936, 287.7471, 
    287.8008, 287.8545, 287.9082, 287.9478, 287.9731, 287.9985, 288.0239, 
    288.0493, 288.0747, 288.0674, 288.0444, 288.0215, 287.9985, 287.9756, 
    287.9526, 287.9299, 287.9158, 287.9016, 287.8877, 287.8735, 287.8596, 
    287.8455, 287.8333, 287.824, 287.8149, 287.8059, 287.7969, 287.7878, 
    287.7769, 287.7642, 287.7512, 287.7385, 287.7256, 287.7129, 287.7, 
    287.6873, 287.6741, 287.6609, 287.6479, 287.6348, 287.6218, 287.6077, 
    287.5935, 287.5796, 287.5654, 287.5515, 287.5374, 287.5232, 287.5093, 
    287.5059, 287.5078, 287.5098, 287.5115, 287.5049, 287.4895, 287.4744, 
    287.459, 287.4438, 287.4285, 287.4131, 287.3979, 287.3826, 287.3586, 
    287.3171, 287.2737, 287.2283, 287.1667, 287.0957, 287.0125, 286.9141, 
    286.7954, 286.6497, 286.467, 286.2305, 284.4067, 284.3315, 284.168, 
    284.0178, 283.8542, 283.668, 283.4817, 283.2954, 283.1091, 282.9231, 
    282.7368, 282.5505, 282.3643, 282.178, 281.9919, 281.8579, 281.7485, 
    281.7744, 281.8003, 281.8262, 281.8521, 281.8779, 281.9038, 281.9297, 
    281.9556, 281.9814, 282.0073, 282.0332, 282.061, 282.0789, 282.0825, 
    282.0862, 282.0896, 282.0933, 282.0969, 282.1003, 282.104, 282.1077, 
    282.1111, 282.1147, 282.1184, 282.1221, 282.1099, 282.0977, 282.0854, 
    282.0732, 282.061, 282.0488, 282.0366, 282.0244, 282.0122, 282, 281.9878, 
    281.9756, 281.9758, 281.9856, 281.9946, 282.0051, 282.0176, 282.032, 
    282.0496, 282.071, 282.0981, 282.1333, 282.1804, 282.2473, 282.3992, 
    282.5388, 282.6699, 282.7944, 282.9189, 283.0435, 283.168, 283.2925, 
    283.417, 283.5415, 283.666, 283.7905, 283.915, 283.9875, 284.0081, 
    284.0281, 284.0186, 284.009, 283.9995, 283.99, 283.9805, 283.9709, 
    283.9614, 283.9519, 283.9424, 283.9329, 283.9287, 283.9246, 283.9204, 
    283.9236, 283.9304, 283.937, 283.9438, 283.9507, 283.9573, 283.9641, 
    283.9707, 283.9775, 283.97, 283.9482, 283.9265, 283.9045, 283.8848, 
    283.8689, 283.8528, 283.8369, 283.8208, 283.8047, 283.7888, 283.7727, 
    283.7568, 283.7393, 283.72, 283.6992, 283.6763, 283.6509, 283.6069, 
    283.5552, 283.4924, 282.2036, 282.1721, 282.1458, 282.1233, 282.0884, 
    282.04, 281.9939, 281.9502, 281.9084, 281.8684, 281.7451, 281.5828, 
    281.4207, 281.2583, 281.0962, 280.9338, 280.7715,
  283.3215, 283.3962, 283.4709, 283.5459, 283.6206, 283.6953, 283.77, 
    283.8447, 283.9197, 283.9944, 284.0691, 284.1138, 284.1433, 284.1445, 
    284.1458, 284.147, 284.1479, 284.1492, 284.1504, 284.1516, 284.1528, 
    284.1541, 284.155, 284.2017, 284.2935, 284.3853, 284.4814, 284.5776, 
    284.6736, 284.7698, 284.866, 284.9622, 285.0581, 285.1543, 285.2505, 
    285.3464, 285.3276, 285.3069, 285.2834, 285.2732, 285.2693, 285.2646, 
    285.259, 285.2522, 285.5862, 285.5867, 285.5872, 285.5876, 285.6416, 
    285.7468, 285.8491, 285.9485, 286.0667, 286.2246, 286.3826, 286.5405, 
    286.6985, 286.8564, 287.0144, 287.1724, 287.3303, 287.3948, 287.4595, 
    287.5242, 287.5889, 287.6533, 287.6973, 287.7412, 287.7854, 287.8293, 
    287.8733, 287.9175, 287.9614, 287.988, 287.9976, 288.0068, 288.0164, 
    288.0256, 288.0349, 288.0242, 288.0039, 287.9834, 287.9631, 287.9429, 
    287.9224, 287.9021, 287.8926, 287.8831, 287.8735, 287.8643, 287.8547, 
    287.8452, 287.8367, 287.8303, 287.824, 287.8174, 287.811, 287.8047, 
    287.7959, 287.7849, 287.7739, 287.7629, 287.752, 287.741, 287.7297, 
    287.7188, 287.7078, 287.6965, 287.6853, 287.6741, 287.6628, 287.6506, 
    287.6382, 287.6257, 287.6135, 287.6011, 287.5886, 287.5762, 287.564, 
    287.5581, 287.5557, 287.553, 287.5505, 287.5374, 287.5137, 287.4902, 
    287.4666, 287.4431, 287.4194, 287.3958, 287.3723, 287.3486, 287.3196, 
    287.2793, 287.238, 287.1953, 287.1338, 287.0627, 286.9797, 286.8821, 
    286.7651, 286.6226, 286.4448, 286.2173, 284.1819, 284.1008, 283.9658, 
    283.8442, 283.7, 283.5237, 283.3474, 283.1709, 282.9946, 282.8184, 
    282.6421, 282.4658, 282.2893, 282.113, 281.9368, 281.7927, 281.6636, 
    281.7004, 281.7371, 281.7739, 281.8108, 281.8474, 281.8843, 281.9209, 
    281.9578, 281.9946, 282.0312, 282.0681, 282.1062, 282.1294, 282.135, 
    282.1409, 282.1467, 282.1523, 282.1582, 282.1638, 282.1697, 282.1753, 
    282.1812, 282.1868, 282.1926, 282.1985, 282.1777, 282.1567, 282.136, 
    282.115, 282.0942, 282.0732, 282.0525, 282.0317, 282.0107, 281.99, 
    281.969, 281.9482, 281.9419, 281.948, 281.9534, 281.9597, 281.967, 
    281.9761, 281.9866, 281.9998, 282.0166, 282.0383, 282.0681, 282.1108, 
    282.1846, 282.3386, 282.4861, 282.6277, 282.7693, 282.9109, 283.0527, 
    283.1943, 283.3359, 283.4775, 283.6194, 283.761, 283.9026, 283.9805, 
    283.9946, 284.0083, 284.0039, 283.9998, 283.9954, 283.991, 283.9866, 
    283.9822, 283.9778, 283.9736, 283.9692, 283.9648, 283.967, 283.9692, 
    283.9714, 283.978, 283.9871, 283.9958, 284.0049, 284.0137, 284.0227, 
    284.0315, 284.0405, 284.0493, 284.0408, 284.0146, 283.9885, 283.9624, 
    283.9375, 283.915, 283.8926, 283.8699, 283.8474, 283.825, 283.8025, 
    283.7798, 283.7573, 283.7324, 283.7051, 283.6743, 283.6399, 283.6006, 
    283.5444, 283.4766, 283.3938, 282.0195, 281.9805, 281.9473, 281.9189, 
    281.8704, 281.8, 281.7319, 281.6658, 281.6013, 281.5388, 281.4221, 
    281.2803, 281.1382, 280.9963, 280.8542, 280.7122, 280.5703,
  283.4966, 283.5537, 283.6111, 283.6682, 283.7256, 283.7827, 283.8398, 
    283.8972, 283.9543, 284.0117, 284.0688, 284.0903, 284.1062, 284.1116, 
    284.1167, 284.1218, 284.1272, 284.1323, 284.1377, 284.1428, 284.1482, 
    284.1533, 284.1584, 284.2175, 284.3301, 284.4426, 284.5566, 284.6709, 
    284.7852, 284.8992, 285.0134, 285.1277, 285.2417, 285.356, 285.4702, 
    285.5842, 285.5769, 285.5686, 285.5591, 285.5557, 285.5557, 285.5554, 
    285.5552, 285.5547, 285.7417, 285.7434, 285.7446, 285.7461, 285.8132, 
    285.9456, 286.0764, 286.2061, 286.3428, 286.4954, 286.6479, 286.8005, 
    286.9531, 287.1057, 287.2583, 287.4109, 287.5635, 287.6057, 287.6477, 
    287.6899, 287.7319, 287.7739, 287.8083, 287.8428, 287.8772, 287.9116, 
    287.9458, 287.9802, 288.0146, 288.0286, 288.022, 288.0151, 288.0085, 
    288.002, 287.9954, 287.9812, 287.9634, 287.9456, 287.9277, 287.9099, 
    287.8921, 287.8743, 287.8694, 287.8645, 287.8596, 287.8547, 287.8499, 
    287.8447, 287.8403, 287.8364, 287.8328, 287.8291, 287.8252, 287.8215, 
    287.8149, 287.8057, 287.7966, 287.7874, 287.7781, 287.7688, 287.7598, 
    287.7505, 287.7412, 287.7319, 287.7227, 287.7134, 287.7041, 287.6934, 
    287.6829, 287.6721, 287.6614, 287.6506, 287.6399, 287.6292, 287.6187, 
    287.6104, 287.6033, 287.5964, 287.5894, 287.5698, 287.5378, 287.5061, 
    287.4741, 287.4424, 287.4104, 287.3784, 287.3467, 287.3147, 287.2808, 
    287.2424, 287.2036, 287.1646, 287.1028, 287.0317, 286.9495, 286.8528, 
    286.7373, 286.5977, 286.4248, 286.2056, 283.9438, 283.8577, 283.7573, 
    283.6692, 283.5457, 283.3794, 283.2129, 283.0466, 282.8801, 282.7136, 
    282.5474, 282.3809, 282.2144, 282.0481, 281.8816, 281.7273, 281.5786, 
    281.6262, 281.6741, 281.7217, 281.7693, 281.8171, 281.8647, 281.9124, 
    281.96, 282.0078, 282.0554, 282.103, 282.1514, 282.1797, 282.1877, 
    282.1956, 282.2036, 282.2114, 282.2195, 282.2273, 282.2351, 282.2432, 
    282.251, 282.259, 282.2668, 282.2749, 282.2454, 282.2158, 282.1863, 
    282.1567, 282.1274, 282.0979, 282.0684, 282.0388, 282.0093, 281.9797, 
    281.9502, 281.9209, 281.9075, 281.9094, 281.9111, 281.9131, 281.9153, 
    281.9182, 281.9214, 281.9255, 281.9307, 281.9377, 281.947, 281.9612, 
    281.9761, 282.1406, 282.3022, 282.4609, 282.6199, 282.7786, 282.9373, 
    283.0962, 283.2549, 283.4138, 283.5725, 283.7312, 283.8901, 283.9734, 
    283.981, 283.9888, 283.9895, 283.9902, 283.9912, 283.9919, 283.9927, 
    283.9937, 283.9944, 283.9951, 283.9961, 283.9968, 284.0054, 284.0139, 
    284.0225, 284.0327, 284.0437, 284.0547, 284.0659, 284.0769, 284.0879, 
    284.0989, 284.1101, 284.1211, 284.1113, 284.0811, 284.0505, 284.0203, 
    283.9902, 283.9612, 283.9321, 283.9031, 283.874, 283.845, 283.8159, 
    283.7869, 283.7578, 283.7256, 283.6892, 283.6477, 283.5999, 283.5439, 
    283.4727, 283.3857, 283.2773, 281.8589, 281.8115, 281.771, 281.7358, 
    281.6726, 281.5784, 281.4851, 281.3926, 281.3013, 281.2109, 281.0991, 
    280.9775, 280.8557, 280.7341, 280.6123, 280.4907, 280.3691,
  283.6189, 283.6597, 283.7007, 283.7415, 283.7825, 283.8232, 283.864, 
    283.905, 283.9458, 283.9868, 284.0276, 284.0413, 284.0552, 284.0688, 
    284.0825, 284.0962, 284.1101, 284.1238, 284.1375, 284.1511, 284.1648, 
    284.1787, 284.1924, 284.2578, 284.376, 284.4946, 284.6145, 284.7351, 
    284.8564, 284.979, 285.1023, 285.2266, 285.3518, 285.4778, 285.605, 
    285.7332, 285.7366, 285.7407, 285.7456, 285.751, 285.7576, 285.7656, 
    285.7751, 285.7874, 285.9258, 285.9282, 285.9304, 285.9324, 286.0049, 
    286.1479, 286.291, 286.4341, 286.5769, 286.72, 286.863, 287.0061, 
    287.1492, 287.2922, 287.4353, 287.5784, 287.7214, 287.7463, 287.7712, 
    287.7961, 287.8213, 287.8462, 287.8711, 287.896, 287.9209, 287.946, 
    287.9709, 287.9958, 288.0208, 288.0264, 288.0127, 287.999, 287.9856, 
    287.9719, 287.9583, 287.9446, 287.9309, 287.9172, 287.9036, 287.8899, 
    287.8762, 287.8625, 287.8601, 287.8577, 287.8555, 287.853, 287.8506, 
    287.8481, 287.8459, 287.8435, 287.8411, 287.8386, 287.8364, 287.834, 
    287.8286, 287.8206, 287.8123, 287.804, 287.7959, 287.7876, 287.7793, 
    287.7712, 287.7629, 287.7549, 287.7466, 287.7383, 287.7302, 287.7205, 
    287.7107, 287.7007, 287.6909, 287.6812, 287.6714, 287.6616, 287.6519, 
    287.6418, 287.6321, 287.6223, 287.6125, 287.5906, 287.5566, 287.5227, 
    287.4885, 287.4546, 287.4207, 287.3865, 287.3525, 287.3186, 287.2847, 
    287.2505, 287.2166, 287.1826, 287.1206, 287.05, 286.9692, 286.8752, 
    286.7654, 286.6345, 286.4766, 286.2815, 283.8411, 283.7485, 283.6692, 
    283.6001, 283.4854, 283.3193, 283.1548, 282.9915, 282.8293, 282.6685, 
    282.5088, 282.3501, 282.1929, 282.0366, 281.8816, 281.7275, 281.5747, 
    281.624, 281.6733, 281.7227, 281.772, 281.8213, 281.8706, 281.9199, 
    281.9692, 282.0183, 282.0676, 282.1169, 282.1663, 282.1968, 282.2085, 
    282.2202, 282.2322, 282.2439, 282.2556, 282.2673, 282.2791, 282.2908, 
    282.3025, 282.3142, 282.3259, 282.3379, 282.302, 282.2661, 282.2302, 
    282.1943, 282.1584, 282.1226, 282.0867, 282.0508, 282.0149, 281.979, 
    281.9431, 281.9072, 281.8916, 281.8967, 281.9028, 281.9099, 281.918, 
    281.9275, 281.939, 281.9529, 281.9702, 281.9927, 282.0225, 282.064, 
    281.8679, 282.041, 282.2131, 282.3838, 282.5532, 282.7212, 282.8882, 
    283.0537, 283.218, 283.3813, 283.5432, 283.7041, 283.8635, 283.9453, 
    283.9497, 283.9543, 283.9587, 283.9634, 283.968, 283.9727, 283.9775, 
    283.9822, 283.9871, 283.9917, 283.9966, 284.0015, 284.0137, 284.0259, 
    284.0381, 284.05, 284.062, 284.0737, 284.0854, 284.0972, 284.1086, 
    284.1201, 284.1316, 284.1428, 284.1326, 284.1006, 284.0684, 284.0359, 
    284.0032, 283.97, 283.9368, 283.9033, 283.8696, 283.8357, 283.8015, 
    283.7671, 283.7322, 283.6929, 283.6477, 283.5955, 283.5347, 283.4624, 
    283.3752, 283.2686, 283.1345, 281.6807, 281.6301, 281.5862, 281.5479, 
    281.479, 281.376, 281.2732, 281.1702, 281.0674, 280.9644, 280.8616, 
    280.7585, 280.6558, 280.5527, 280.45, 280.3469, 280.2441,
  283.6621, 283.6885, 283.7148, 283.741, 283.7673, 283.7937, 283.8198, 
    283.8462, 283.8726, 283.8987, 283.925, 283.9539, 283.9829, 284.0117, 
    284.0405, 284.0696, 284.0984, 284.1272, 284.1562, 284.1851, 284.2139, 
    284.2429, 284.2717, 284.3357, 284.4368, 284.5405, 284.6472, 284.7566, 
    284.8689, 284.9846, 285.1033, 285.2256, 285.3513, 285.4807, 285.614, 
    286.0127, 286.0444, 286.0691, 286.0889, 286.1052, 286.1187, 286.1299, 
    286.1399, 286.1482, 286.1558, 286.1621, 286.168, 286.1733, 286.2393, 
    286.3665, 286.4937, 286.6211, 286.7483, 286.8755, 287.0027, 287.1299, 
    287.2571, 287.3845, 287.5117, 287.6389, 287.7661, 287.782, 287.7979, 
    287.8137, 287.8296, 287.8455, 287.8613, 287.8772, 287.8931, 287.9089, 
    287.9248, 287.9407, 287.9565, 287.9607, 287.9536, 287.9463, 287.9392, 
    287.9321, 287.9248, 287.9177, 287.9104, 287.9033, 287.896, 287.8889, 
    287.8816, 287.8745, 287.8716, 287.8687, 287.866, 287.863, 287.8601, 
    287.8572, 287.8545, 287.8516, 287.8486, 287.8457, 287.8428, 287.8401, 
    287.8345, 287.8259, 287.8176, 287.8091, 287.8008, 287.7922, 287.7839, 
    287.7756, 287.7671, 287.7588, 287.7502, 287.7419, 287.7336, 287.7234, 
    287.7134, 287.7031, 287.6931, 287.6831, 287.6729, 287.6628, 287.6528, 
    287.6426, 287.6326, 287.6226, 287.6123, 287.594, 287.5671, 287.5403, 
    287.5134, 287.4866, 287.4597, 287.4329, 287.406, 287.3792, 287.3523, 
    287.3254, 287.2986, 287.2717, 287.208, 287.137, 287.0574, 286.9673, 
    286.865, 286.7476, 286.6113, 286.4514, 286.261, 286.0308, 285.7463, 
    285.3862, 285.0889, 284.9224, 284.7432, 284.5493, 282.8792, 282.7163, 
    282.5579, 282.4038, 282.2539, 282.1079, 281.9658, 281.8271, 281.6924, 
    281.7292, 281.7664, 281.8032, 281.8403, 281.8772, 281.9143, 281.9514, 
    281.9883, 282.0254, 282.0623, 282.0994, 282.1362, 282.1638, 282.1819, 
    282.2, 282.218, 282.2361, 282.2542, 282.2722, 282.2903, 282.3083, 
    282.3264, 282.3445, 282.3625, 282.3806, 282.3418, 282.3027, 282.2639, 
    282.2251, 282.186, 282.1472, 282.1084, 282.0693, 282.0305, 281.9917, 
    281.9529, 281.9138, 281.9033, 281.9229, 281.9446, 281.9692, 281.9968, 
    282.0286, 282.0652, 282.1079, 282.1582, 282.2188, 282.2925, 282.385, 
    282.5037, 282.5671, 282.6357, 282.7097, 282.7898, 282.8767, 282.9717, 
    283.0754, 283.1895, 283.3965, 283.54, 283.6797, 283.8159, 283.8853, 
    283.8904, 283.8958, 283.9014, 283.907, 283.9128, 283.9189, 283.925, 
    283.9314, 283.9377, 283.9446, 283.9514, 283.3445, 283.3792, 283.4165, 
    283.4565, 283.5, 283.5474, 283.5989, 283.6553, 283.7173, 284.0605, 
    284.0706, 284.0801, 284.0894, 284.0791, 284.0488, 284.0178, 283.9858, 
    283.3203, 283.1931, 283.0774, 282.9714, 282.8745, 282.7852, 282.7026, 
    282.6262, 282.5552, 282.313, 282.1248, 281.9741, 281.8508, 281.748, 
    281.6609, 281.5864, 281.5217, 281.4651, 281.4153, 281.3708, 281.3311, 
    281.2695, 281.1833, 281.0969, 281.0105, 280.9241, 280.8379, 280.7515, 
    280.665, 280.5786, 280.4922, 280.406, 280.3196, 280.2332,
  283.7053, 283.717, 283.7288, 283.7405, 283.7522, 283.7639, 283.7756, 
    283.7874, 283.7991, 283.8108, 283.8225, 283.8667, 283.9106, 283.9546, 
    283.9988, 284.0427, 284.0869, 284.1309, 284.175, 284.219, 284.2629, 
    284.3071, 284.3511, 284.4143, 284.4995, 284.5889, 284.6821, 284.78, 
    284.8828, 284.991, 285.1045, 285.2244, 285.3506, 285.4841, 285.6255, 
    286.0991, 286.1484, 286.1907, 286.2266, 286.2581, 286.2856, 286.3098, 
    286.3315, 286.3508, 286.3684, 286.3843, 286.3987, 286.4119, 286.4736, 
    286.5852, 286.6965, 286.8079, 286.9194, 287.0308, 287.1423, 287.2537, 
    287.3652, 287.4766, 287.5879, 287.6995, 287.8108, 287.8176, 287.8245, 
    287.8311, 287.8379, 287.8447, 287.8516, 287.8582, 287.865, 287.8718, 
    287.8784, 287.8853, 287.8921, 287.895, 287.8943, 287.8936, 287.8928, 
    287.8921, 287.8916, 287.8909, 287.8901, 287.8894, 287.8887, 287.8879, 
    287.8872, 287.8865, 287.8831, 287.8796, 287.8765, 287.873, 287.8696, 
    287.8662, 287.8628, 287.8596, 287.8562, 287.8528, 287.8494, 287.8462, 
    287.8401, 287.8315, 287.823, 287.8142, 287.8057, 287.7971, 287.7886, 
    287.7798, 287.7712, 287.7627, 287.7542, 287.7454, 287.7368, 287.7266, 
    287.7161, 287.7058, 287.6953, 287.6851, 287.6746, 287.6643, 287.6538, 
    287.6433, 287.6331, 287.6226, 287.6123, 287.5972, 287.5776, 287.5579, 
    287.5381, 287.5186, 287.4988, 287.479, 287.4595, 287.4397, 287.4199, 
    287.4004, 287.3806, 287.3608, 287.2937, 287.2205, 287.1399, 287.0513, 
    286.9531, 286.844, 286.7219, 286.584, 286.4277, 286.2483, 286.041, 
    285.7983, 285.594, 285.4507, 285.2927, 285.1172, 282.9377, 282.7712, 
    282.613, 282.4629, 282.3198, 282.1833, 282.0532, 281.9287, 281.8098, 
    281.8345, 281.8594, 281.884, 281.9087, 281.9333, 281.958, 281.9829, 
    282.0076, 282.0322, 282.0569, 282.0815, 282.1064, 282.1309, 282.1553, 
    282.1797, 282.2041, 282.2283, 282.2527, 282.2771, 282.3015, 282.3259, 
    282.3503, 282.3745, 282.3989, 282.4233, 282.3816, 282.3396, 282.2976, 
    282.2559, 282.2139, 282.1721, 282.1301, 282.0881, 282.0464, 282.0044, 
    281.9626, 281.9207, 281.9153, 281.9482, 281.9844, 282.0242, 282.0679, 
    282.1165, 282.1709, 282.2317, 282.3008, 282.3794, 282.47, 282.5754, 
    282.6997, 282.7395, 282.7832, 282.8318, 282.886, 282.9465, 283.0146, 
    283.0923, 283.1814, 283.4128, 283.5366, 283.6548, 283.7678, 283.8247, 
    283.8296, 283.8347, 283.8398, 283.8455, 283.8513, 283.8574, 283.864, 
    283.8708, 283.8779, 283.8855, 283.8936, 283.1421, 283.1738, 283.209, 
    283.2478, 283.291, 283.3394, 283.3938, 283.4558, 283.5271, 284.0093, 
    284.0183, 284.0271, 284.0354, 284.0251, 283.9958, 283.9648, 283.9326, 
    282.9846, 282.8381, 282.7104, 282.5981, 282.4985, 282.4097, 282.3298, 
    282.2576, 282.1921, 282.0217, 281.8772, 281.7532, 281.6453, 281.5505, 
    281.467, 281.3926, 281.3259, 281.2656, 281.2112, 281.1616, 281.1165, 
    281.0603, 280.9905, 280.9207, 280.8508, 280.781, 280.7112, 280.6414, 
    280.5715, 280.5017, 280.4319, 280.3621, 280.2922, 280.2224,
  283.7488, 283.7458, 283.7429, 283.7402, 283.7373, 283.7344, 283.7314, 
    283.7285, 283.7258, 283.7229, 283.72, 283.7793, 283.8384, 283.8977, 
    283.9568, 284.0161, 284.0752, 284.1345, 284.1936, 284.2529, 284.3123, 
    284.3713, 284.4307, 284.4937, 284.5642, 284.6394, 284.7197, 284.8059, 
    284.8984, 284.998, 285.106, 285.2229, 285.3499, 285.4888, 285.6409, 
    286.1519, 286.2175, 286.2764, 286.3296, 286.3782, 286.4221, 286.4626, 
    286.4998, 286.5342, 286.5657, 286.5952, 286.6226, 286.6482, 286.708, 
    286.8037, 286.8994, 286.9949, 287.0906, 287.1863, 287.2817, 287.3774, 
    287.4731, 287.5686, 287.6643, 287.76, 287.8557, 287.8533, 287.8508, 
    287.8486, 287.8462, 287.844, 287.8416, 287.8394, 287.8369, 287.8347, 
    287.8323, 287.8301, 287.8276, 287.8293, 287.8352, 287.8408, 287.8467, 
    287.8523, 287.8582, 287.864, 287.8696, 287.8755, 287.8811, 287.887, 
    287.8926, 287.8984, 287.8945, 287.8906, 287.8867, 287.8831, 287.8792, 
    287.8752, 287.8713, 287.8677, 287.8638, 287.8599, 287.856, 287.8523, 
    287.8459, 287.8372, 287.8281, 287.8193, 287.8105, 287.8018, 287.793, 
    287.7842, 287.7754, 287.7666, 287.7578, 287.749, 287.7402, 287.7295, 
    287.7188, 287.7083, 287.6975, 287.6868, 287.6763, 287.6655, 287.6548, 
    287.644, 287.6335, 287.6228, 287.6121, 287.6006, 287.5881, 287.5754, 
    287.563, 287.5503, 287.5378, 287.5254, 287.5127, 287.5002, 287.4878, 
    287.4751, 287.4626, 287.4502, 287.3779, 287.3005, 287.2175, 287.1282, 
    287.0317, 286.9272, 286.814, 286.6904, 286.5554, 286.4067, 286.2429, 
    286.061, 285.906, 285.7834, 285.6458, 285.4905, 283.0076, 282.8352, 
    282.6758, 282.5283, 282.3911, 282.2634, 282.144, 282.0322, 281.9275, 
    281.9397, 281.9521, 281.9646, 281.9771, 281.9895, 282.002, 282.0144, 
    282.0266, 282.0391, 282.0515, 282.064, 282.0764, 282.0979, 282.1287, 
    282.1592, 282.1899, 282.2207, 282.2515, 282.282, 282.3127, 282.3435, 
    282.374, 282.4048, 282.4355, 282.4661, 282.4214, 282.3765, 282.3315, 
    282.2866, 282.2417, 282.1968, 282.1519, 282.1069, 282.0623, 282.0173, 
    281.9724, 281.9275, 281.9268, 281.9729, 282.022, 282.075, 282.1321, 
    282.1936, 282.2605, 282.3333, 282.4126, 282.4998, 282.5955, 282.7017, 
    282.8196, 282.8467, 282.877, 282.9111, 282.95, 282.9941, 283.0452, 
    283.1047, 283.175, 283.4304, 283.5332, 283.6292, 283.7192, 283.7637, 
    283.7668, 283.7705, 283.7742, 283.7781, 283.7825, 283.7871, 283.7922, 
    283.7976, 283.8035, 283.8098, 283.8169, 283.0181, 283.0459, 283.0769, 
    283.1118, 283.1516, 283.197, 283.2493, 283.3105, 283.3828, 283.9541, 
    283.9639, 283.9727, 283.981, 283.9709, 283.9412, 283.9094, 283.8755, 
    282.73, 282.5793, 282.4519, 282.3428, 282.2483, 282.1655, 282.0925, 
    282.0278, 281.9697, 281.8289, 281.7021, 281.5879, 281.4839, 281.3892, 
    281.3022, 281.2224, 281.1487, 281.0806, 281.0173, 280.9585, 280.9038, 
    280.8511, 280.7976, 280.7444, 280.6912, 280.6379, 280.5845, 280.5312, 
    280.478, 280.4246, 280.3713, 280.3181, 280.2649, 280.2114,
  283.792, 283.7747, 283.7571, 283.7397, 283.7222, 283.7048, 283.6873, 
    283.6699, 283.6523, 283.635, 283.6174, 283.6919, 283.7661, 283.8406, 
    283.915, 283.9893, 284.0637, 284.1382, 284.2124, 284.2869, 284.3613, 
    284.4355, 284.51, 284.5737, 284.6306, 284.6924, 284.76, 284.8342, 
    284.916, 285.0066, 285.1077, 285.2209, 285.3489, 285.4946, 285.6621, 
    286.1875, 286.2664, 286.3403, 286.4097, 286.4749, 286.5361, 286.594, 
    286.6487, 286.7004, 286.7495, 286.7959, 286.8401, 286.8823, 286.9424, 
    287.0222, 287.1021, 287.1819, 287.2617, 287.3416, 287.4214, 287.5012, 
    287.5811, 287.6609, 287.7407, 287.8206, 287.9004, 287.8889, 287.8774, 
    287.866, 287.8547, 287.8433, 287.8318, 287.8203, 287.8091, 287.7976, 
    287.7861, 287.7747, 287.7634, 287.7637, 287.7759, 287.7881, 287.8003, 
    287.8125, 287.8247, 287.8369, 287.8494, 287.8616, 287.8738, 287.886, 
    287.8982, 287.9104, 287.906, 287.9016, 287.8972, 287.8931, 287.8887, 
    287.8843, 287.8799, 287.8757, 287.8713, 287.8669, 287.8625, 287.8582, 
    287.8516, 287.8425, 287.8335, 287.8245, 287.8157, 287.8066, 287.7976, 
    287.7886, 287.7795, 287.7705, 287.7615, 287.7524, 287.7434, 287.7327, 
    287.7217, 287.7107, 287.6997, 287.6887, 287.6777, 287.6667, 287.6558, 
    287.6448, 287.634, 287.623, 287.6121, 287.6038, 287.5984, 287.593, 
    287.5876, 287.5823, 287.5769, 287.5715, 287.5662, 287.5608, 287.5554, 
    287.55, 287.5447, 287.5393, 287.4604, 287.3777, 287.2905, 287.1987, 
    287.1021, 287, 286.8921, 286.7776, 286.6562, 286.5273, 286.3899, 
    286.2434, 286.1179, 286.012, 285.8918, 285.7546, 283.0925, 282.9104, 
    282.7476, 282.6013, 282.4688, 282.3484, 282.2383, 282.1377, 282.0449, 
    282.0452, 282.0452, 282.0454, 282.0454, 282.0457, 282.0457, 282.0459, 
    282.0459, 282.0461, 282.0461, 282.0461, 282.0464, 282.0649, 282.1021, 
    282.1389, 282.176, 282.2129, 282.25, 282.2869, 282.324, 282.3608, 
    282.3979, 282.4351, 282.4719, 282.509, 282.4612, 282.4131, 282.3652, 
    282.3174, 282.2695, 282.2217, 282.1738, 282.1257, 282.0779, 282.03, 
    281.9822, 281.9343, 281.9385, 281.9966, 282.0579, 282.1223, 282.1904, 
    282.262, 282.3376, 282.418, 282.5029, 282.593, 282.689, 282.7913, 
    282.9006, 282.9202, 282.9419, 282.9668, 282.9956, 283.0288, 283.0676, 
    283.114, 283.1704, 283.4492, 283.5293, 283.6028, 283.6702, 283.7019, 
    283.7024, 283.7029, 283.7034, 283.7041, 283.7046, 283.7053, 283.7063, 
    283.707, 283.7083, 283.7092, 283.7107, 282.9343, 282.9583, 282.9856, 
    283.0166, 283.0522, 283.0935, 283.1418, 283.1997, 283.2695, 283.895, 
    283.9062, 283.9167, 283.926, 283.916, 283.885, 283.8511, 283.814, 
    282.5303, 282.3821, 282.2598, 282.1572, 282.0696, 281.9941, 281.9285, 
    281.8708, 281.8198, 281.6917, 281.572, 281.4595, 281.354, 281.2544, 
    281.1606, 281.0718, 280.988, 280.9084, 280.833, 280.7612, 280.6929, 
    280.6416, 280.605, 280.5681, 280.5315, 280.4946, 280.458, 280.4211, 
    280.3845, 280.3477, 280.311, 280.2742, 280.2375, 280.2007,
  283.8352, 283.8032, 283.7712, 283.7393, 283.7073, 283.675, 283.6431, 
    283.6111, 283.5791, 283.5469, 283.5149, 283.6045, 283.6941, 283.7834, 
    283.873, 283.9626, 284.0522, 284.1416, 284.2312, 284.3208, 284.4104, 
    284.4998, 284.5894, 284.6545, 284.699, 284.7483, 284.8032, 284.8655, 
    284.9358, 285.0166, 285.1096, 285.2188, 285.3477, 285.5029, 285.6934, 
    286.2131, 286.303, 286.3896, 286.4734, 286.5544, 286.6326, 286.708, 
    286.7812, 286.8521, 286.9207, 286.9873, 287.0518, 287.1143, 287.177, 
    287.241, 287.3049, 287.3689, 287.4329, 287.4971, 287.561, 287.625, 
    287.689, 287.7529, 287.8171, 287.8811, 287.9451, 287.9246, 287.9041, 
    287.8835, 287.863, 287.8425, 287.822, 287.8015, 287.781, 287.7605, 
    287.74, 287.7195, 287.699, 287.698, 287.7168, 287.7354, 287.7542, 
    287.7727, 287.7915, 287.8101, 287.8289, 287.8477, 287.8662, 287.885, 
    287.9036, 287.9224, 287.9175, 287.9126, 287.9077, 287.9031, 287.8982, 
    287.8933, 287.8884, 287.8835, 287.8789, 287.874, 287.8691, 287.8643, 
    287.8574, 287.8481, 287.8389, 287.8296, 287.8206, 287.8113, 287.802, 
    287.793, 287.7837, 287.7744, 287.7654, 287.7561, 287.7468, 287.7356, 
    287.7244, 287.7131, 287.7019, 287.6907, 287.6794, 287.6682, 287.657, 
    287.6455, 287.6343, 287.623, 287.6118, 287.6072, 287.6089, 287.6106, 
    287.6125, 287.6143, 287.616, 287.6179, 287.6196, 287.6213, 287.6233, 
    287.625, 287.6267, 287.6287, 287.5415, 287.4519, 287.3594, 287.2639, 
    287.1655, 287.064, 286.959, 286.8503, 286.7383, 286.6221, 286.5017, 
    286.3772, 286.2712, 286.1787, 286.0732, 285.9514, 283.1978, 283.0005, 
    282.8306, 282.6829, 282.5535, 282.4387, 282.3367, 282.2451, 282.1626, 
    282.1504, 282.1382, 282.126, 282.1138, 282.1016, 282.0894, 282.0774, 
    282.0652, 282.053, 282.0408, 282.0286, 282.0164, 282.032, 282.0752, 
    282.1187, 282.1619, 282.2053, 282.2485, 282.2917, 282.3352, 282.3784, 
    282.4219, 282.4651, 282.5085, 282.5518, 282.501, 282.45, 282.3992, 
    282.3481, 282.2974, 282.2463, 282.1956, 282.1445, 282.0938, 282.0427, 
    281.9919, 281.9409, 281.9497, 282.02, 282.092, 282.1667, 282.2434, 
    282.3228, 282.4048, 282.4895, 282.5769, 282.6675, 282.7612, 282.8584, 
    282.959, 282.9734, 282.9895, 283.0083, 283.0298, 283.0552, 283.0852, 
    283.1216, 283.1665, 283.4695, 283.5254, 283.5757, 283.6206, 283.6396, 
    283.636, 283.6318, 283.6274, 283.6221, 283.6162, 283.6096, 283.6018, 
    283.5925, 283.5818, 283.5688, 283.553, 282.8738, 282.8948, 282.9187, 
    282.946, 282.9778, 283.0149, 283.0591, 283.1125, 283.1785, 283.8313, 
    283.8459, 283.8589, 283.8706, 283.8606, 283.8269, 283.7898, 283.748, 
    282.3691, 282.2268, 282.1116, 282.0161, 281.9358, 281.8674, 281.8083, 
    281.7568, 281.7117, 281.5891, 281.4712, 281.3572, 281.2468, 281.1404, 
    281.0374, 280.9377, 280.8413, 280.7478, 280.6572, 280.5693, 280.4841, 
    280.4324, 280.4121, 280.3918, 280.3718, 280.3516, 280.3313, 280.311, 
    280.291, 280.2708, 280.2505, 280.2302, 280.21, 280.1899,
  283.8787, 283.832, 283.7854, 283.7388, 283.6921, 283.6455, 283.5989, 
    283.5522, 283.5056, 283.459, 283.4124, 283.5171, 283.6218, 283.7266, 
    283.8311, 283.9358, 284.0405, 284.1453, 284.25, 284.3547, 284.4595, 
    284.564, 284.6687, 284.7363, 284.7693, 284.8071, 284.8501, 284.9001, 
    284.9587, 285.0283, 285.1123, 285.2156, 285.3459, 285.5154, 285.7449, 
    286.2327, 286.3315, 286.4292, 286.5256, 286.6208, 286.7151, 286.8081, 
    286.9001, 286.991, 287.0808, 287.1697, 287.2576, 287.3442, 287.4114, 
    287.4595, 287.5078, 287.5559, 287.6042, 287.6523, 287.7007, 287.7488, 
    287.7969, 287.8452, 287.8933, 287.9417, 287.9897, 287.9602, 287.9307, 
    287.9011, 287.8713, 287.8418, 287.8123, 287.7827, 287.7529, 287.7234, 
    287.6938, 287.6643, 287.6345, 287.6323, 287.6575, 287.6826, 287.7078, 
    287.7329, 287.7581, 287.7832, 287.8083, 287.8335, 287.8589, 287.884, 
    287.9092, 287.9343, 287.929, 287.9236, 287.9182, 287.9131, 287.9077, 
    287.9023, 287.897, 287.8916, 287.8865, 287.8811, 287.8757, 287.8704, 
    287.863, 287.8538, 287.8442, 287.835, 287.8254, 287.8159, 287.8066, 
    287.7971, 287.7878, 287.7783, 287.769, 287.7595, 287.7502, 287.7388, 
    287.7271, 287.7156, 287.7041, 287.6926, 287.6809, 287.6694, 287.658, 
    287.6462, 287.6348, 287.6233, 287.6118, 287.6104, 287.6194, 287.6284, 
    287.6372, 287.6462, 287.6553, 287.6641, 287.6731, 287.6819, 287.6909, 
    287.7, 287.7087, 287.7178, 287.6211, 287.5234, 287.4243, 287.3245, 
    287.2231, 287.1206, 287.0171, 286.9121, 286.8059, 286.6985, 286.5898, 
    286.4797, 286.3872, 286.3059, 286.2124, 286.1038, 283.3318, 283.1096, 
    282.9275, 282.7751, 282.646, 282.5352, 282.439, 282.3545, 282.28, 
    282.2556, 282.2312, 282.2065, 282.1821, 282.1577, 282.1333, 282.1086, 
    282.0842, 282.0598, 282.0354, 282.011, 281.9863, 281.999, 282.0486, 
    282.0981, 282.1479, 282.1975, 282.2471, 282.2969, 282.3464, 282.396, 
    282.4456, 282.4954, 282.5449, 282.5945, 282.5408, 282.4868, 282.4329, 
    282.3789, 282.325, 282.2712, 282.2173, 282.1633, 282.1094, 282.0557, 
    282.0017, 281.9478, 281.9612, 282.0425, 282.1248, 282.208, 282.2922, 
    282.3774, 282.4636, 282.5508, 282.6392, 282.7285, 282.8188, 282.9104, 
    283.0032, 283.0139, 283.0259, 283.04, 283.0564, 283.0757, 283.0991, 
    283.1274, 283.1633, 283.4912, 283.5212, 283.5476, 283.5706, 283.5769, 
    283.5676, 283.5571, 283.5452, 283.5312, 283.5149, 283.4954, 283.4719, 
    283.4431, 283.4067, 283.3594, 283.2952, 282.8284, 282.8467, 282.8674, 
    282.8916, 282.9197, 282.9531, 282.9932, 283.042, 283.1033, 283.7627, 
    283.7825, 283.7996, 283.8147, 283.8047, 283.7673, 283.7251, 283.6765, 
    282.2368, 282.1016, 281.9934, 281.9053, 281.8318, 281.7695, 281.7163, 
    281.6702, 281.6299, 281.5098, 281.3909, 281.2734, 281.1575, 281.0427, 
    280.9294, 280.8176, 280.707, 280.5977, 280.4895, 280.3828, 280.2771, 
    280.2231, 280.2195, 280.2158, 280.2119, 280.2083, 280.2046, 280.2009, 
    280.1973, 280.1936, 280.1899, 280.1863, 280.1826, 280.179,
  283.8945, 283.8474, 283.8005, 283.7534, 283.7065, 283.6594, 283.6125, 
    283.5657, 283.5186, 283.4717, 283.4246, 283.5298, 283.6357, 283.7422, 
    283.8496, 283.9578, 284.0664, 284.176, 284.2864, 284.3975, 284.5095, 
    284.6221, 284.7356, 284.8057, 284.835, 284.8684, 284.9072, 284.9531, 
    285.0078, 285.0742, 285.1567, 285.262, 285.4004, 285.5913, 285.8706, 
    286.3196, 286.418, 286.5164, 286.6147, 286.7131, 286.8115, 286.9099, 
    287.0083, 287.1067, 287.2051, 287.3035, 287.4019, 287.5002, 287.5679, 
    287.6042, 287.6406, 287.6772, 287.7136, 287.7502, 287.7866, 287.823, 
    287.8596, 287.896, 287.9326, 287.969, 288.0056, 287.9712, 287.937, 
    287.9028, 287.8687, 287.8345, 287.8003, 287.7661, 287.7319, 287.6978, 
    287.6636, 287.6294, 287.5952, 287.592, 287.6204, 287.6484, 287.6765, 
    287.7046, 287.7327, 287.761, 287.7891, 287.8171, 287.8452, 287.8733, 
    287.9016, 287.9297, 287.9241, 287.9185, 287.9126, 287.907, 287.9014, 
    287.8958, 287.8901, 287.8845, 287.8789, 287.873, 287.8674, 287.8618, 
    287.8547, 287.8462, 287.8374, 287.8289, 287.8203, 287.8118, 287.803, 
    287.7944, 287.7859, 287.7773, 287.7686, 287.76, 287.7515, 287.7397, 
    287.728, 287.7166, 287.7048, 287.6931, 287.6814, 287.6699, 287.6582, 
    287.6465, 287.6348, 287.6233, 287.6116, 287.6123, 287.6255, 287.6389, 
    287.6521, 287.6653, 287.6785, 287.6917, 287.7051, 287.7183, 287.7314, 
    287.7446, 287.7581, 287.7712, 287.6716, 287.572, 287.4724, 287.3728, 
    287.2732, 287.1736, 287.074, 286.9744, 286.8748, 286.7751, 286.6755, 
    286.5759, 286.4922, 286.4172, 286.3308, 286.2302, 283.5002, 283.2566, 
    283.0637, 282.907, 282.7773, 282.6682, 282.575, 282.4946, 282.4246, 
    282.3875, 282.3506, 282.3137, 282.2766, 282.2397, 282.2029, 282.166, 
    282.1289, 282.092, 282.0552, 282.0181, 281.9812, 281.989, 282.0417, 
    282.0942, 282.147, 282.1995, 282.252, 282.3047, 282.3572, 282.4099, 
    282.4624, 282.5149, 282.5676, 282.6201, 282.5696, 282.5193, 282.4688, 
    282.4182, 282.3677, 282.3171, 282.2666, 282.2161, 282.1655, 282.1152, 
    282.0647, 282.0142, 282.0317, 282.1172, 282.2026, 282.2883, 282.3738, 
    282.4592, 282.5449, 282.6304, 282.7158, 282.8015, 282.887, 282.9724, 
    283.0579, 283.0645, 283.0718, 283.0801, 283.0898, 283.1013, 283.115, 
    283.1313, 283.1516, 283.4988, 283.5107, 283.5212, 283.5303, 283.5273, 
    283.512, 283.4939, 283.4731, 283.4487, 283.4194, 283.3838, 283.3396, 
    283.2834, 283.2095, 283.1074, 282.9578, 282.7178, 282.7273, 282.7383, 
    282.751, 282.7654, 282.7825, 282.803, 282.8276, 282.8579, 283.6787, 
    283.7053, 283.728, 283.7478, 283.7373, 283.6943, 283.6448, 283.5872, 
    282.0054, 281.895, 281.8059, 281.7322, 281.6704, 281.6177, 281.5723, 
    281.5325, 281.4978, 281.3816, 281.2651, 281.1489, 281.0325, 280.9163, 
    280.8, 280.6836, 280.5674, 280.4509, 280.3347, 280.2185, 280.1021, 
    280.0469, 280.053, 280.0588, 280.0649, 280.071, 280.0769, 280.083, 
    280.0889, 280.095, 280.1008, 280.1069, 280.1128, 280.1189,
  283.864, 283.8408, 283.8174, 283.7939, 283.7708, 283.7473, 283.7239, 
    283.7007, 283.6772, 283.6538, 283.6306, 283.7136, 283.7988, 283.8862, 
    283.9761, 284.0684, 284.1628, 284.26, 284.3601, 284.4629, 284.5686, 
    284.6772, 284.7891, 284.8628, 284.8989, 284.9404, 284.9883, 285.0439, 
    285.1101, 285.1897, 285.2871, 285.4092, 285.5667, 285.7778, 286.0757, 
    286.5266, 286.6106, 286.6946, 286.7786, 286.8625, 286.9465, 287.0308, 
    287.1147, 287.1987, 287.2827, 287.3667, 287.4507, 287.5347, 287.5925, 
    287.6243, 287.6558, 287.6875, 287.719, 287.7507, 287.7825, 287.814, 
    287.8457, 287.8772, 287.9089, 287.9404, 287.9722, 287.9409, 287.9097, 
    287.8787, 287.8474, 287.8162, 287.7849, 287.7539, 287.7227, 287.6914, 
    287.6602, 287.6289, 287.5979, 287.5947, 287.6201, 287.6453, 287.6704, 
    287.6956, 287.7207, 287.7461, 287.7712, 287.7964, 287.8215, 287.8467, 
    287.8718, 287.8972, 287.8914, 287.8857, 287.8799, 287.8743, 287.8687, 
    287.8628, 287.8572, 287.8513, 287.8457, 287.8401, 287.8342, 287.8286, 
    287.8225, 287.8164, 287.8103, 287.8042, 287.7981, 287.792, 287.7859, 
    287.7798, 287.7737, 287.7676, 287.7615, 287.7554, 287.7493, 287.7378, 
    287.7263, 287.7148, 287.7031, 287.6917, 287.6802, 287.6687, 287.6572, 
    287.6458, 287.6343, 287.6228, 287.6111, 287.6118, 287.6245, 287.6372, 
    287.6499, 287.6626, 287.6753, 287.688, 287.7007, 287.7134, 287.7261, 
    287.7388, 287.7515, 287.7642, 287.675, 287.5857, 287.4963, 287.407, 
    287.3179, 287.2285, 287.1392, 287.05, 286.9607, 286.8713, 286.7822, 
    286.6929, 286.6147, 286.541, 286.4561, 286.3572, 283.6724, 283.4326, 
    283.2429, 283.0889, 282.9612, 282.854, 282.7622, 282.6831, 282.6143, 
    282.5645, 282.5149, 282.4651, 282.4155, 282.3657, 282.3162, 282.2664, 
    282.2168, 282.167, 282.1172, 282.0676, 282.0178, 282.0181, 282.0679, 
    282.1179, 282.1677, 282.2175, 282.2676, 282.3174, 282.3674, 282.4172, 
    282.467, 282.5171, 282.5669, 282.6169, 282.5806, 282.5442, 282.5078, 
    282.4717, 282.4353, 282.3989, 282.3625, 282.3262, 282.29, 282.2537, 
    282.2173, 282.1809, 282.2021, 282.2808, 282.3591, 282.4377, 282.5164, 
    282.5947, 282.6733, 282.752, 282.8306, 282.9089, 282.9875, 283.0662, 
    283.1448, 283.1436, 283.1423, 283.1409, 283.1392, 283.1375, 283.1353, 
    283.1328, 283.1299, 283.4758, 283.4861, 283.4951, 283.5029, 283.4963, 
    283.4744, 283.4492, 283.4202, 283.386, 283.3457, 283.2974, 283.238, 
    283.1638, 283.0676, 282.9392, 282.7578, 282.4832, 282.4768, 282.4697, 
    282.4619, 282.4529, 282.4426, 282.4309, 282.4172, 282.4011, 283.5603, 
    283.5938, 283.6226, 283.6479, 283.636, 283.5842, 283.5249, 283.4565, 
    281.6489, 281.5718, 281.5063, 281.4497, 281.4006, 281.3574, 281.3193, 
    281.2852, 281.2546, 281.1482, 281.042, 280.9355, 280.8291, 280.7229, 
    280.6165, 280.51, 280.4038, 280.2974, 280.1909, 280.0847, 279.9783, 
    279.927, 279.9312, 279.9351, 279.9392, 279.9431, 279.9473, 279.9512, 
    279.9553, 279.9592, 279.9634, 279.9675, 279.9714, 279.9756,
  283.8337, 283.834, 283.8342, 283.8345, 283.8347, 283.835, 283.8354, 
    283.8357, 283.8359, 283.8362, 283.8364, 283.9009, 283.9683, 284.0388, 
    284.1128, 284.1902, 284.2715, 284.3569, 284.4468, 285.5833, 285.6768, 
    285.7607, 285.8369, 285.9426, 286.0662, 286.1714, 286.2625, 286.3416, 
    286.4114, 286.4731, 286.5281, 286.5776, 286.6223, 286.6628, 286.6997, 
    286.7336, 286.8032, 286.8728, 286.9424, 287.0122, 287.0818, 287.1514, 
    287.2209, 287.2905, 287.3604, 287.4299, 287.4995, 287.5691, 287.6174, 
    287.6443, 287.6709, 287.6978, 287.7246, 287.7512, 287.7781, 287.8049, 
    287.8318, 287.8584, 287.8853, 287.9121, 287.9387, 287.9106, 287.8823, 
    287.8542, 287.8259, 287.7979, 287.7698, 287.7415, 287.7134, 287.6851, 
    287.657, 287.6287, 287.6006, 287.5974, 287.6199, 287.6421, 287.6643, 
    287.6865, 287.7087, 287.731, 287.7534, 287.7756, 287.7979, 287.8201, 
    287.8423, 287.8645, 287.8589, 287.853, 287.8472, 287.8416, 287.8357, 
    287.8298, 287.8242, 287.8184, 287.8125, 287.8069, 287.801, 287.7952, 
    287.7905, 287.7869, 287.7832, 287.7795, 287.7761, 287.7725, 287.7688, 
    287.7651, 287.7615, 287.7578, 287.7542, 287.7507, 287.7471, 287.7356, 
    287.7244, 287.7129, 287.7017, 287.6902, 287.679, 287.6675, 287.6562, 
    287.6448, 287.6335, 287.6221, 287.6108, 287.6113, 287.6233, 287.6355, 
    287.6477, 287.6599, 287.6721, 287.6843, 287.6965, 287.7085, 287.7207, 
    287.7329, 287.7451, 287.7573, 287.6782, 287.5994, 287.5203, 287.4414, 
    287.3625, 287.2834, 287.2046, 287.1255, 287.0466, 286.9675, 286.8887, 
    286.8096, 286.7373, 286.6648, 286.5813, 286.4839, 283.8442, 283.6089, 
    283.4221, 283.2708, 283.1453, 283.0396, 282.9497, 282.8718, 282.804, 
    282.7417, 282.6792, 282.6167, 282.5542, 282.4917, 282.4292, 282.3669, 
    282.3044, 282.2419, 282.1794, 282.1169, 282.0547, 282.0469, 282.0942, 
    282.1414, 282.1887, 282.2358, 282.283, 282.3303, 282.3774, 282.4246, 
    282.4719, 282.519, 282.5664, 282.6135, 282.5913, 282.5693, 282.5471, 
    282.5249, 282.5029, 282.4807, 282.4585, 282.4365, 282.4143, 282.3921, 
    282.3701, 282.3479, 282.3726, 282.4441, 282.5156, 282.5872, 282.6589, 
    282.7305, 282.802, 282.8735, 282.9451, 283.0166, 283.0881, 283.1599, 
    283.2314, 283.2212, 283.21, 283.1978, 283.1843, 283.1692, 283.1526, 
    283.134, 283.1128, 283.0889, 283.0615, 283.0295, 282.9922, 282.9124, 
    282.8086, 282.7202, 282.644, 282.5776, 282.519, 282.4673, 282.4211, 
    282.3796, 282.342, 282.3081, 282.2771, 282.2488, 282.2312, 282.2119, 
    282.1909, 282.1677, 282.1421, 282.1135, 282.0813, 282.0452, 282.0039, 
    281.9568, 281.9021, 281.8379, 281.7373, 281.6238, 281.5271, 281.4438, 
    281.3711, 281.3071, 281.2505, 281.2, 281.1545, 281.1135, 281.0764, 
    281.0425, 281.0115, 280.915, 280.8186, 280.7222, 280.6257, 280.5293, 
    280.4329, 280.3364, 280.24, 280.1436, 280.0471, 279.9507, 279.8542, 
    279.8071, 279.8093, 279.8113, 279.8135, 279.8154, 279.8176, 279.8196, 
    279.8218, 279.8237, 279.8259, 279.8279, 279.8301, 279.832,
  283.8032, 283.8271, 283.8511, 283.875, 283.8989, 283.9229, 283.9468, 
    283.9707, 283.9946, 284.0183, 284.0422, 284.0918, 284.1443, 284.2004, 
    284.2607, 284.3252, 284.3945, 284.4692, 284.55, 285.7971, 285.874, 
    285.9421, 286.0029, 286.0916, 286.2031, 286.3037, 286.3945, 286.4773, 
    286.5527, 286.6221, 286.6858, 286.7446, 286.7991, 286.8496, 286.8967, 
    286.9407, 286.9958, 287.051, 287.1064, 287.1616, 287.2168, 287.2722, 
    287.3274, 287.3826, 287.4377, 287.4932, 287.5483, 287.6035, 287.6421, 
    287.6641, 287.686, 287.708, 287.73, 287.752, 287.7739, 287.7957, 
    287.8176, 287.8396, 287.8616, 287.8835, 287.9055, 287.8804, 287.855, 
    287.8298, 287.8047, 287.7795, 287.7544, 287.729, 287.7039, 287.6787, 
    287.6536, 287.6284, 287.6033, 287.6003, 287.6196, 287.6389, 287.6582, 
    287.6775, 287.6968, 287.7161, 287.7356, 287.7549, 287.7742, 287.7935, 
    287.8127, 287.832, 287.8262, 287.8203, 287.8145, 287.8086, 287.803, 
    287.7971, 287.7913, 287.7854, 287.7795, 287.7737, 287.7678, 287.762, 
    287.7583, 287.7573, 287.7561, 287.7551, 287.7539, 287.7527, 287.7517, 
    287.7505, 287.7493, 287.7483, 287.7471, 287.7458, 287.7449, 287.7336, 
    287.7224, 287.7112, 287.7, 287.6887, 287.6777, 287.6665, 287.6553, 
    287.644, 287.6328, 287.6216, 287.6104, 287.6106, 287.6223, 287.634, 
    287.6455, 287.6572, 287.6689, 287.6804, 287.6921, 287.7039, 287.7153, 
    287.7271, 287.7388, 287.7502, 287.6816, 287.613, 287.5444, 287.4758, 
    287.407, 287.3384, 287.2698, 287.2012, 287.1326, 287.0637, 286.9951, 
    286.9265, 286.8599, 286.7886, 286.7065, 286.6108, 284.0164, 283.7849, 
    283.6013, 283.4524, 283.3291, 283.2253, 283.137, 283.0605, 282.9939, 
    282.9187, 282.8435, 282.7683, 282.6929, 282.6177, 282.5425, 282.4673, 
    282.3921, 282.3169, 282.2417, 282.1665, 282.0913, 282.0759, 282.1204, 
    282.165, 282.2095, 282.2539, 282.2986, 282.343, 282.3875, 282.4321, 
    282.4766, 282.5212, 282.5657, 282.6101, 282.6023, 282.5942, 282.5864, 
    282.5784, 282.5703, 282.5625, 282.5544, 282.5466, 282.5386, 282.5305, 
    282.5227, 282.5146, 282.543, 282.6077, 282.6721, 282.7368, 282.8013, 
    282.866, 282.9307, 282.9951, 283.0598, 283.1243, 283.189, 283.2534, 
    283.3181, 283.2974, 283.2751, 283.2512, 283.2256, 283.1978, 283.1677, 
    283.135, 283.0994, 283.0603, 283.0173, 282.9697, 282.917, 282.8303, 
    282.7229, 282.6262, 282.5388, 282.4595, 282.387, 282.3203, 282.259, 
    282.2026, 282.1501, 282.1016, 282.0564, 282.0142, 281.99, 281.9641, 
    281.9365, 281.9065, 281.8743, 281.8394, 281.8013, 281.7598, 281.7144, 
    281.6646, 281.6094, 281.5481, 281.4651, 281.3733, 281.291, 281.2163, 
    281.1484, 281.0864, 281.0298, 280.9775, 280.9292, 280.8845, 280.843, 
    280.8044, 280.7683, 280.6819, 280.5955, 280.5088, 280.4224, 280.3359, 
    280.2493, 280.1628, 280.0764, 279.99, 279.9033, 279.8169, 279.7305, 
    279.6873, 279.6873, 279.6875, 279.6875, 279.6877, 279.6877, 279.688, 
    279.688, 279.6882, 279.6882, 279.6885, 279.6885, 279.6887,
  283.7729, 283.8203, 283.8679, 283.9155, 283.9631, 284.0105, 284.0581, 
    284.1057, 284.1531, 284.2007, 284.2483, 284.2861, 284.3274, 284.3723, 
    284.4214, 284.4756, 284.5352, 284.6016, 284.6755, 285.948, 286.0112, 
    286.0664, 286.1152, 286.1946, 286.3027, 286.4041, 286.499, 286.5884, 
    286.6726, 286.752, 286.8269, 286.8979, 286.9653, 287.0291, 287.0898, 
    287.1477, 287.1885, 287.2292, 287.2703, 287.311, 287.3521, 287.3928, 
    287.4336, 287.4746, 287.5154, 287.5564, 287.5972, 287.6379, 287.667, 
    287.6841, 287.7012, 287.7183, 287.7354, 287.7524, 287.7695, 287.7866, 
    287.8037, 287.8208, 287.8379, 287.855, 287.8721, 287.8499, 287.8276, 
    287.8057, 287.7834, 287.7612, 287.739, 287.7168, 287.6946, 287.6724, 
    287.6501, 287.6279, 287.6057, 287.603, 287.6194, 287.6357, 287.6521, 
    287.6685, 287.6848, 287.7012, 287.7175, 287.7341, 287.7505, 287.7668, 
    287.7832, 287.7996, 287.7937, 287.7878, 287.7817, 287.7759, 287.77, 
    287.7642, 287.7583, 287.7522, 287.7463, 287.7405, 287.7346, 287.7285, 
    287.7263, 287.7278, 287.729, 287.7305, 287.7317, 287.7332, 287.7344, 
    287.7358, 287.7371, 287.7385, 287.7397, 287.7412, 287.7427, 287.7314, 
    287.7205, 287.7095, 287.6985, 287.6873, 287.6763, 287.6653, 287.6543, 
    287.6433, 287.6321, 287.6211, 287.6101, 287.6101, 287.6213, 287.6323, 
    287.6436, 287.6545, 287.6658, 287.6768, 287.688, 287.699, 287.7102, 
    287.7212, 287.7322, 287.7434, 287.6851, 287.6267, 287.5684, 287.51, 
    287.4517, 287.3933, 287.335, 287.2766, 287.2183, 287.1599, 287.1016, 
    287.0432, 286.9824, 286.9124, 286.8318, 286.7378, 284.1885, 283.9609, 
    283.7805, 283.6343, 283.5132, 283.4111, 283.3242, 283.249, 283.1836, 
    283.0957, 283.0076, 282.9197, 282.8318, 282.7437, 282.6558, 282.5679, 
    282.4797, 282.3918, 282.304, 282.2158, 282.1279, 282.1047, 282.1467, 
    282.1885, 282.2305, 282.2722, 282.314, 282.356, 282.3977, 282.4395, 
    282.4814, 282.5232, 282.5649, 282.6069, 282.613, 282.6194, 282.6255, 
    282.6318, 282.6379, 282.6443, 282.6504, 282.6567, 282.6628, 282.6692, 
    282.6753, 282.6816, 282.7136, 282.771, 282.8286, 282.8862, 282.9438, 
    283.0015, 283.0591, 283.1167, 283.1743, 283.2319, 283.2896, 283.3472, 
    283.4048, 283.3721, 283.3376, 283.3015, 283.2634, 283.2231, 283.1807, 
    283.1357, 283.0881, 283.0376, 282.9836, 282.9263, 282.865, 282.7734, 
    282.6606, 282.5549, 282.4558, 282.3625, 282.2749, 282.1921, 282.114, 
    282.04, 281.9697, 281.9031, 281.8398, 281.7795, 281.7534, 281.7258, 
    281.697, 281.6665, 281.6343, 281.6001, 281.5642, 281.5259, 281.4854, 
    281.4424, 281.3965, 281.3474, 281.2766, 281.1914, 281.1113, 281.0364, 
    280.9661, 280.8997, 280.8372, 280.7781, 280.7219, 280.6689, 280.6187, 
    280.5708, 280.5251, 280.4487, 280.3721, 280.2954, 280.219, 280.1423, 
    280.0659, 279.9893, 279.9128, 279.8362, 279.7595, 279.6831, 279.6064, 
    279.5674, 279.5654, 279.5637, 279.5618, 279.5601, 279.5581, 279.5564, 
    279.5544, 279.5527, 279.5508, 279.5491, 279.5471, 279.5454,
  283.7424, 283.8137, 283.8848, 283.9561, 284.0271, 284.0984, 284.1694, 
    284.2407, 284.3118, 284.3831, 284.4541, 284.4844, 284.5178, 284.5549, 
    284.5967, 284.644, 284.6978, 284.7593, 284.8311, 286.0603, 286.1123, 
    286.1572, 286.1965, 286.27, 286.3784, 286.4829, 286.5837, 286.6812, 
    286.7754, 286.8662, 286.9543, 287.0396, 287.1221, 287.2019, 287.2795, 
    287.3547, 287.3811, 287.4077, 287.4341, 287.4607, 287.4871, 287.5137, 
    287.54, 287.5664, 287.593, 287.6194, 287.646, 287.6724, 287.6919, 
    287.7041, 287.7163, 287.7285, 287.7407, 287.7529, 287.7654, 287.7776, 
    287.7898, 287.802, 287.8142, 287.8264, 287.8389, 287.8196, 287.8003, 
    287.7812, 287.762, 287.7429, 287.7236, 287.7043, 287.6853, 287.666, 
    287.647, 287.6277, 287.6084, 287.6057, 287.6191, 287.6326, 287.646, 
    287.6594, 287.6729, 287.6863, 287.6997, 287.7134, 287.7268, 287.7402, 
    287.7537, 287.7671, 287.761, 287.7551, 287.749, 287.7432, 287.7371, 
    287.7312, 287.7251, 287.7192, 287.7131, 287.7073, 287.7012, 287.6953, 
    287.6943, 287.698, 287.7019, 287.7058, 287.7095, 287.7134, 287.7173, 
    287.7212, 287.7249, 287.7288, 287.7327, 287.7366, 287.7402, 287.7295, 
    287.7185, 287.7078, 287.6968, 287.686, 287.675, 287.6641, 287.6533, 
    287.6423, 287.6316, 287.6206, 287.6099, 287.6096, 287.6201, 287.6309, 
    287.6414, 287.6519, 287.6624, 287.6731, 287.6836, 287.6941, 287.7048, 
    287.7153, 287.7258, 287.7366, 287.6885, 287.6404, 287.5923, 287.5444, 
    287.4963, 287.4482, 287.4004, 287.3523, 287.3042, 287.2561, 287.2083, 
    287.1602, 287.105, 287.0361, 286.957, 286.8645, 284.3604, 284.137, 
    283.9597, 283.8162, 283.697, 283.5969, 283.5115, 283.4377, 283.3735, 
    283.2727, 283.1719, 283.0713, 282.9705, 282.8699, 282.769, 282.6682, 
    282.5676, 282.4668, 282.366, 282.2654, 282.1646, 282.1338, 282.1729, 
    282.2122, 282.2512, 282.2903, 282.3296, 282.3687, 282.4077, 282.447, 
    282.4861, 282.5251, 282.5645, 282.6035, 282.624, 282.6443, 282.6648, 
    282.6851, 282.7056, 282.7261, 282.7463, 282.7668, 282.7871, 282.8076, 
    282.8281, 282.8484, 282.884, 282.9346, 282.9851, 283.0359, 283.0864, 
    283.1372, 283.1877, 283.2383, 283.2891, 283.3396, 283.3901, 283.4409, 
    283.4915, 283.4453, 283.3979, 283.3489, 283.2983, 283.2461, 283.1921, 
    283.1365, 283.0789, 283.019, 282.9573, 282.8933, 282.8269, 282.7317, 
    282.6133, 282.4988, 282.3884, 282.282, 282.179, 282.0793, 281.9832, 
    281.8899, 281.7996, 281.7122, 281.6274, 281.5452, 281.5212, 281.4966, 
    281.4712, 281.4448, 281.4177, 281.3899, 281.3608, 281.3308, 281.3, 
    281.2678, 281.2346, 281.2002, 281.1384, 281.053, 280.9705, 280.8906, 
    280.8137, 280.7395, 280.6677, 280.5981, 280.5308, 280.4656, 280.4026, 
    280.3413, 280.282, 280.2153, 280.1487, 280.0823, 280.0156, 279.949, 
    279.8823, 279.8157, 279.749, 279.6824, 279.616, 279.5493, 279.4827, 
    279.4475, 279.4436, 279.4399, 279.436, 279.4321, 279.4285, 279.4246, 
    279.4209, 279.417, 279.4133, 279.4094, 279.4058, 279.4019,
  283.7122, 283.8069, 283.9016, 283.9966, 284.0913, 284.186, 284.2808, 
    284.3757, 284.4705, 284.5652, 284.6602, 284.6863, 284.7161, 284.7498, 
    284.7888, 284.834, 284.8875, 284.9512, 285.0288, 286.1472, 286.1897, 
    286.2261, 286.2578, 286.3279, 286.4377, 286.5466, 286.6538, 286.7598, 
    286.8643, 286.9678, 287.0698, 287.1707, 287.27, 287.3684, 287.4656, 
    287.5618, 287.5737, 287.5859, 287.5979, 287.6101, 287.6221, 287.6343, 
    287.6465, 287.6584, 287.6707, 287.6826, 287.6948, 287.7068, 287.7166, 
    287.7241, 287.7314, 287.7388, 287.7463, 287.7537, 287.761, 287.7683, 
    287.7759, 287.7832, 287.7905, 287.7981, 287.8054, 287.7893, 287.7729, 
    287.7568, 287.7407, 287.7244, 287.7083, 287.6921, 287.676, 287.6597, 
    287.6436, 287.6274, 287.6111, 287.6084, 287.6189, 287.6294, 287.6399, 
    287.6504, 287.6609, 287.6714, 287.6819, 287.6924, 287.7031, 287.7136, 
    287.7241, 287.7346, 287.7285, 287.7224, 287.7163, 287.7104, 287.7043, 
    287.6982, 287.6921, 287.6863, 287.6802, 287.6741, 287.668, 287.6619, 
    287.6621, 287.6685, 287.6748, 287.6812, 287.6875, 287.6938, 287.7002, 
    287.7065, 287.7129, 287.7192, 287.7253, 287.7317, 287.738, 287.7273, 
    287.7166, 287.7061, 287.6953, 287.6846, 287.6738, 287.6631, 287.6523, 
    287.6416, 287.6309, 287.6201, 287.6094, 287.6091, 287.6191, 287.6292, 
    287.6392, 287.6492, 287.6592, 287.6692, 287.6792, 287.6895, 287.6995, 
    287.7095, 287.7195, 287.7295, 287.6919, 287.6541, 287.6165, 287.5786, 
    287.541, 287.5032, 287.4656, 287.4277, 287.3901, 287.3523, 287.3147, 
    287.2771, 287.2275, 287.1602, 287.0823, 286.9915, 284.5325, 284.313, 
    284.1392, 283.998, 283.8811, 283.7827, 283.6987, 283.6265, 283.5632, 
    283.4497, 283.3362, 283.2227, 283.1091, 282.9958, 282.8823, 282.7688, 
    282.6553, 282.5417, 282.4282, 282.3147, 282.2012, 282.1628, 282.1992, 
    282.2356, 282.2722, 282.3086, 282.345, 282.3813, 282.418, 282.4543, 
    282.4907, 282.5273, 282.5637, 282.6001, 282.6348, 282.6694, 282.7039, 
    282.7385, 282.7732, 282.8079, 282.8423, 282.877, 282.9116, 282.946, 
    282.9807, 283.0154, 283.0544, 283.0981, 283.1418, 283.1853, 283.229, 
    283.2727, 283.3164, 283.3599, 283.4036, 283.4473, 283.491, 283.5344, 
    283.5781, 283.5173, 283.4561, 283.3938, 283.3308, 283.2671, 283.2024, 
    283.137, 283.0708, 283.0039, 282.936, 282.8672, 282.7976, 282.7, 
    282.5759, 282.4536, 282.3328, 282.2136, 282.0957, 281.9795, 281.8645, 
    281.751, 281.6389, 281.5281, 281.4187, 281.3105, 281.2932, 281.2756, 
    281.2578, 281.24, 281.2217, 281.2034, 281.1846, 281.1658, 281.1465, 
    281.1272, 281.1077, 281.0876, 281.033, 280.9443, 280.8567, 280.7703, 
    280.6848, 280.6006, 280.5173, 280.4353, 280.354, 280.2737, 280.1946, 
    280.1162, 280.0388, 279.9822, 279.9255, 279.8689, 279.8123, 279.7554, 
    279.6987, 279.6421, 279.5854, 279.5288, 279.4722, 279.4153, 279.3586, 
    279.3274, 279.3218, 279.3159, 279.3103, 279.3044, 279.2988, 279.293, 
    279.2874, 279.2815, 279.2759, 279.27, 279.2642, 279.2585,
  283.75, 283.8528, 283.9563, 284.0605, 284.1655, 284.271, 284.3772, 
    284.4841, 284.5918, 284.7002, 284.8091, 284.8369, 284.8687, 284.9053, 
    284.9482, 284.999, 285.0603, 285.1355, 285.23, 286.2573, 286.2942, 
    286.3264, 286.3545, 286.4207, 286.5276, 286.6345, 286.7415, 286.8484, 
    286.9553, 287.0623, 287.1692, 287.2764, 287.3833, 287.4902, 287.5972, 
    287.7041, 287.7065, 287.7092, 287.7117, 287.7144, 287.7168, 287.7195, 
    287.7219, 287.7246, 287.7273, 287.7297, 287.7324, 287.7349, 287.739, 
    287.7446, 287.7502, 287.7559, 287.7615, 287.7671, 287.7727, 287.7783, 
    287.7839, 287.7896, 287.7949, 287.8005, 287.8062, 287.791, 287.7759, 
    287.7605, 287.7454, 287.7302, 287.7148, 287.6997, 287.6846, 287.6692, 
    287.6541, 287.6389, 287.6235, 287.6194, 287.626, 287.6326, 287.6394, 
    287.646, 287.6526, 287.6592, 287.666, 287.6726, 287.6792, 287.6858, 
    287.6926, 287.6992, 287.6943, 287.6897, 287.6848, 287.6799, 287.6753, 
    287.6704, 287.6658, 287.6609, 287.656, 287.6514, 287.6465, 287.6418, 
    287.6433, 287.6511, 287.6589, 287.6667, 287.6746, 287.6821, 287.6899, 
    287.6978, 287.7056, 287.7134, 287.7212, 287.729, 287.7368, 287.7268, 
    287.7166, 287.7063, 287.6963, 287.686, 287.676, 287.6658, 287.6558, 
    287.6455, 287.6353, 287.6252, 287.615, 287.6143, 287.623, 287.6316, 
    287.6404, 287.6489, 287.6577, 287.6663, 287.675, 287.6836, 287.6924, 
    287.7009, 287.7097, 287.7183, 287.6897, 287.6609, 287.6321, 287.6035, 
    287.5747, 287.5459, 287.5173, 287.4885, 287.4597, 287.4312, 287.4023, 
    287.3735, 287.3301, 287.2656, 287.1914, 287.105, 284.76, 284.5508, 
    284.385, 284.2505, 284.1389, 284.0452, 283.9651, 283.896, 283.8359, 
    283.7065, 283.5774, 283.448, 283.3188, 283.1895, 283.0603, 282.9309, 
    282.8018, 282.6724, 282.5432, 282.4138, 282.2847, 282.2346, 282.2639, 
    282.2935, 282.3228, 282.3521, 282.3813, 282.4109, 282.4402, 282.4695, 
    282.499, 282.5283, 282.5576, 282.5869, 282.6292, 282.6714, 282.7136, 
    282.7559, 282.7979, 282.8401, 282.8823, 282.9246, 282.9668, 283.0088, 
    283.051, 283.0933, 283.1333, 283.1709, 283.2085, 283.2463, 283.2839, 
    283.3218, 283.3594, 283.397, 283.4348, 283.4724, 283.5103, 283.5479, 
    283.5854, 283.5156, 283.4456, 283.3757, 283.3057, 283.2358, 283.1658, 
    283.0959, 283.0259, 282.9561, 282.886, 282.8162, 282.7461, 282.6494, 
    282.5261, 282.4028, 282.2793, 282.156, 282.0325, 281.9092, 281.7859, 
    281.6624, 281.5391, 281.4158, 281.2922, 281.1689, 281.1543, 281.1399, 
    281.1255, 281.1108, 281.0964, 281.0818, 281.0674, 281.0527, 281.0383, 
    281.0239, 281.0093, 280.9949, 280.9424, 280.8523, 280.762, 280.6719, 
    280.5815, 280.4915, 280.4011, 280.311, 280.2207, 280.1306, 280.0403, 
    279.9502, 279.8599, 279.8115, 279.7629, 279.7146, 279.666, 279.6177, 
    279.5691, 279.5208, 279.4724, 279.4238, 279.3755, 279.3269, 279.2786, 
    279.25, 279.2415, 279.2327, 279.2241, 279.2156, 279.2068, 279.1982, 
    279.1897, 279.1809, 279.1724, 279.1638, 279.1553, 279.1465,
  283.9236, 284.0061, 284.0908, 284.178, 284.2671, 284.3589, 284.4531, 
    284.5498, 284.6494, 284.7517, 284.8569, 284.8911, 284.9302, 284.9749, 
    285.0266, 285.0879, 285.1606, 285.249, 285.3586, 286.4309, 286.4712, 
    286.5068, 286.5388, 286.6003, 286.6938, 286.7874, 286.8811, 286.9746, 
    287.0681, 287.1616, 287.2551, 287.3489, 287.4424, 287.5359, 287.6294, 
    287.7229, 287.7253, 287.7275, 287.73, 287.7322, 287.7344, 287.7368, 
    287.739, 287.7415, 287.7437, 287.7458, 287.7483, 287.7505, 287.7566, 
    287.7661, 287.7759, 287.7854, 287.7952, 287.8049, 287.8145, 287.8242, 
    287.8337, 287.8435, 287.853, 287.8628, 287.8723, 287.8542, 287.8362, 
    287.8181, 287.7998, 287.7817, 287.7637, 287.7454, 287.7273, 287.7092, 
    287.6912, 287.6729, 287.6548, 287.6462, 287.6472, 287.6482, 287.6492, 
    287.6504, 287.6514, 287.6523, 287.6533, 287.6543, 287.6553, 287.6562, 
    287.6572, 287.6584, 287.6575, 287.6565, 287.6553, 287.6543, 287.6533, 
    287.6523, 287.6514, 287.6504, 287.6494, 287.6484, 287.6475, 287.6465, 
    287.6497, 287.657, 287.6643, 287.6716, 287.679, 287.6863, 287.6936, 
    287.7009, 287.7083, 287.7156, 287.7229, 287.73, 287.7373, 287.7285, 
    287.72, 287.7112, 287.7024, 287.6936, 287.6848, 287.676, 287.6672, 
    287.6584, 287.6497, 287.6409, 287.6321, 287.6306, 287.6362, 287.6421, 
    287.6477, 287.6536, 287.6592, 287.6648, 287.6707, 287.6763, 287.6821, 
    287.6877, 287.6934, 287.6992, 287.6768, 287.6545, 287.6323, 287.6099, 
    287.5876, 287.5654, 287.543, 287.5208, 287.4985, 287.4761, 287.4539, 
    287.4314, 287.3943, 287.3367, 287.2703, 287.1929, 285.094, 284.9067, 
    284.7583, 284.6379, 284.5381, 284.4541, 284.3826, 284.3208, 284.2668, 
    284.116, 283.9653, 283.8145, 283.6636, 283.5127, 283.3621, 283.2112, 
    283.0603, 282.9094, 282.7588, 282.6079, 282.457, 282.3887, 282.4026, 
    282.4163, 282.4302, 282.4441, 282.458, 282.4719, 282.4856, 282.4995, 
    282.5134, 282.5273, 282.5413, 282.5552, 282.5923, 282.6294, 282.6665, 
    282.7039, 282.741, 282.7781, 282.8154, 282.8525, 282.8896, 282.927, 
    282.9641, 283.0012, 283.0366, 283.0706, 283.1042, 283.1379, 283.1716, 
    283.2053, 283.239, 283.2727, 283.3064, 283.3401, 283.374, 283.4077, 
    283.4414, 283.3748, 283.3081, 283.2415, 283.1748, 283.1082, 283.0417, 
    282.9751, 282.9084, 282.8418, 282.7751, 282.7085, 282.6421, 282.5525, 
    282.4402, 282.3279, 282.2156, 282.1033, 281.991, 281.8787, 281.7664, 
    281.6541, 281.5417, 281.4294, 281.3171, 281.2048, 281.1794, 281.1541, 
    281.1287, 281.1033, 281.0779, 281.0525, 281.0273, 281.002, 280.9766, 
    280.9512, 280.9258, 280.9004, 280.8445, 280.7576, 280.6709, 280.5842, 
    280.4973, 280.4106, 280.324, 280.2373, 280.1504, 280.0637, 279.9771, 
    279.8901, 279.8035, 279.76, 279.7166, 279.6731, 279.6296, 279.5862, 
    279.5427, 279.4993, 279.4558, 279.4124, 279.3689, 279.3254, 279.282, 
    279.2534, 279.2402, 279.2271, 279.2139, 279.2004, 279.1873, 279.1741, 
    279.1609, 279.1475, 279.1343, 279.1211, 279.1079, 279.0945,
  284.1055, 284.1699, 284.2375, 284.3083, 284.3828, 284.4609, 284.5432, 
    284.6296, 284.7212, 284.8176, 284.9197, 284.9619, 285.0098, 285.0642, 
    285.127, 285.2, 285.2859, 285.3889, 285.5142, 286.5916, 286.6389, 
    286.6821, 286.7217, 286.78, 286.8604, 286.9404, 287.0205, 287.1006, 
    287.1809, 287.261, 287.3411, 287.4214, 287.5015, 287.5815, 287.6616, 
    287.7419, 287.7439, 287.7458, 287.748, 287.75, 287.752, 287.7542, 
    287.7561, 287.7581, 287.7603, 287.7622, 287.7642, 287.7664, 287.7742, 
    287.7878, 287.8015, 287.8152, 287.8289, 287.8425, 287.8564, 287.8701, 
    287.8838, 287.8975, 287.9111, 287.9248, 287.9385, 287.9175, 287.8965, 
    287.8755, 287.8542, 287.8333, 287.8123, 287.7913, 287.7703, 287.749, 
    287.728, 287.707, 287.686, 287.6731, 287.6685, 287.6638, 287.6592, 
    287.6545, 287.6499, 287.6453, 287.6406, 287.636, 287.6313, 287.6267, 
    287.6221, 287.6174, 287.6204, 287.623, 287.626, 287.6287, 287.6316, 
    287.6343, 287.6372, 287.6401, 287.6428, 287.6458, 287.6484, 287.6514, 
    287.656, 287.6628, 287.6697, 287.6765, 287.6833, 287.6902, 287.697, 
    287.7039, 287.7107, 287.7175, 287.7244, 287.7312, 287.738, 287.7305, 
    287.7231, 287.7158, 287.7085, 287.7009, 287.6936, 287.6863, 287.6787, 
    287.6714, 287.6641, 287.6567, 287.6492, 287.647, 287.6497, 287.6523, 
    287.6553, 287.658, 287.6606, 287.6636, 287.6663, 287.6689, 287.6716, 
    287.6746, 287.6772, 287.6799, 287.6641, 287.6482, 287.6323, 287.6165, 
    287.6006, 287.5847, 287.5688, 287.553, 287.5371, 287.5212, 287.5054, 
    287.4895, 287.4585, 287.4077, 287.3489, 287.2805, 285.428, 285.2627, 
    285.1316, 285.0254, 284.9373, 284.8633, 284.8, 284.7454, 284.698, 
    284.5256, 284.3533, 284.1809, 284.0085, 283.8362, 283.6638, 283.4915, 
    283.3191, 283.1467, 282.9744, 282.802, 282.6296, 282.5425, 282.541, 
    282.5393, 282.5378, 282.5361, 282.5344, 282.533, 282.5312, 282.5295, 
    282.5281, 282.5264, 282.5247, 282.5232, 282.5552, 282.5874, 282.6196, 
    282.6519, 282.6841, 282.7163, 282.7483, 282.7805, 282.8127, 282.845, 
    282.8772, 282.9094, 282.9402, 282.97, 282.9998, 283.0295, 283.0593, 
    283.0889, 283.1187, 283.1484, 283.1782, 283.208, 283.2375, 283.2673, 
    283.2971, 283.2339, 283.1707, 283.1072, 283.0439, 282.9807, 282.9175, 
    282.8542, 282.7908, 282.7275, 282.6643, 282.6011, 282.5378, 282.4556, 
    282.3542, 282.2529, 282.1519, 282.0505, 281.9492, 281.8481, 281.7468, 
    281.6455, 281.5444, 281.4431, 281.3418, 281.2405, 281.2043, 281.1682, 
    281.1321, 281.0957, 281.0596, 281.0234, 280.9871, 280.9509, 280.9148, 
    280.8787, 280.8423, 280.8062, 280.7463, 280.6631, 280.5798, 280.4966, 
    280.4133, 280.3301, 280.2468, 280.1633, 280.0801, 279.9968, 279.9136, 
    279.8303, 279.7471, 279.7085, 279.6702, 279.6316, 279.593, 279.5547, 
    279.5161, 279.4775, 279.4392, 279.4006, 279.3621, 279.3237, 279.2852, 
    279.2571, 279.2393, 279.2212, 279.2034, 279.1855, 279.1677, 279.1499, 
    279.1318, 279.114, 279.0962, 279.0784, 279.0605, 279.0427,
  284.2964, 284.3455, 284.3982, 284.4546, 284.5154, 284.5811, 284.6521, 
    284.729, 284.813, 284.9048, 285.0056, 285.0581, 285.1169, 285.1833, 
    285.259, 285.3457, 285.4465, 285.5649, 285.7061, 286.7405, 286.7986, 
    286.8525, 286.9026, 286.96, 287.0266, 287.0933, 287.1602, 287.2268, 
    287.2937, 287.3604, 287.427, 287.4939, 287.5605, 287.6272, 287.6941, 
    287.7607, 287.7625, 287.7644, 287.7661, 287.7678, 287.7695, 287.7715, 
    287.7732, 287.7749, 287.7766, 287.7783, 287.7803, 287.782, 287.7917, 
    287.8096, 287.8271, 287.845, 287.8628, 287.8804, 287.8982, 287.916, 
    287.9336, 287.9514, 287.9692, 287.9868, 288.0046, 287.9807, 287.9568, 
    287.9329, 287.9089, 287.885, 287.8608, 287.8369, 287.813, 287.7891, 
    287.7651, 287.7412, 287.7173, 287.7002, 287.6897, 287.6794, 287.6692, 
    287.6589, 287.6487, 287.6384, 287.6282, 287.6177, 287.6074, 287.5972, 
    287.5869, 287.5767, 287.5833, 287.5898, 287.5964, 287.603, 287.6096, 
    287.6165, 287.623, 287.6296, 287.6362, 287.6428, 287.6494, 287.656, 
    287.6626, 287.6689, 287.6753, 287.6816, 287.6877, 287.6941, 287.7004, 
    287.7068, 287.7131, 287.7195, 287.7258, 287.7322, 287.7385, 287.7324, 
    287.7266, 287.7205, 287.7144, 287.7085, 287.7024, 287.6963, 287.6904, 
    287.6843, 287.6785, 287.6724, 287.6663, 287.6633, 287.6631, 287.6628, 
    287.6626, 287.6624, 287.6621, 287.6621, 287.6619, 287.6616, 287.6614, 
    287.6611, 287.6611, 287.6609, 287.6514, 287.6418, 287.6326, 287.623, 
    287.6135, 287.604, 287.5947, 287.5852, 287.5757, 287.5662, 287.5569, 
    287.5474, 287.5227, 287.4785, 287.4277, 287.3684, 285.762, 285.6187, 
    285.5051, 285.4128, 285.3364, 285.2722, 285.2175, 285.1702, 285.1289, 
    284.9351, 284.7412, 284.5471, 284.3533, 284.1594, 283.9656, 283.7715, 
    283.5776, 283.3838, 283.1899, 282.9961, 282.802, 282.6965, 282.6794, 
    282.6624, 282.6453, 282.6282, 282.6111, 282.5938, 282.5767, 282.5596, 
    282.5425, 282.5254, 282.5083, 282.4912, 282.5183, 282.5454, 282.5728, 
    282.5999, 282.627, 282.6543, 282.6814, 282.7085, 282.7358, 282.7629, 
    282.79, 282.8174, 282.8438, 282.8696, 282.8953, 282.9211, 282.9468, 
    282.9727, 282.9983, 283.0242, 283.0498, 283.0757, 283.1013, 283.1272, 
    283.1528, 283.093, 283.033, 282.9731, 282.9131, 282.8533, 282.7932, 
    282.7334, 282.6733, 282.6133, 282.5535, 282.4934, 282.4336, 282.3584, 
    282.2683, 282.1782, 282.0879, 281.9978, 281.9077, 281.8174, 281.7273, 
    281.6372, 281.5469, 281.4568, 281.3667, 281.2764, 281.2295, 281.1824, 
    281.1353, 281.0881, 281.0413, 280.9941, 280.947, 280.8999, 280.853, 
    280.8059, 280.7588, 280.7119, 280.6484, 280.5686, 280.4888, 280.4089, 
    280.3291, 280.2493, 280.1694, 280.0896, 280.0098, 279.9302, 279.8503, 
    279.7705, 279.6907, 279.6572, 279.6235, 279.5901, 279.5566, 279.5232, 
    279.4895, 279.4561, 279.4226, 279.3892, 279.3555, 279.322, 279.2886, 
    279.2605, 279.238, 279.2156, 279.1931, 279.1707, 279.1482, 279.1255, 
    279.103, 279.0806, 279.0581, 279.0356, 279.0132, 278.9907,
  284.4971, 284.5342, 285.4729, 285.5854, 285.6785, 285.7566, 285.8232, 
    285.8806, 285.9307, 285.9749, 286.0137, 286.136, 286.2505, 286.3574, 
    286.4578, 286.5522, 286.6411, 286.7249, 286.8042, 286.8792, 286.9504, 
    287.0178, 287.082, 287.1396, 287.1929, 287.2463, 287.2996, 287.353, 
    287.4062, 287.4597, 287.5129, 287.5664, 287.6196, 287.6731, 287.7263, 
    287.7798, 287.7812, 287.7827, 287.7842, 287.7856, 287.7871, 287.7886, 
    287.79, 287.7917, 287.7932, 287.7947, 287.7961, 287.7976, 287.8093, 
    287.8311, 287.8528, 287.8748, 287.8965, 287.9182, 287.9399, 287.9619, 
    287.9836, 288.0054, 288.0271, 288.0491, 288.0708, 288.0439, 288.0171, 
    287.9902, 287.9634, 287.9365, 287.9097, 287.8828, 287.856, 287.8291, 
    287.802, 287.7751, 287.7483, 287.7271, 287.7109, 287.6951, 287.6792, 
    287.6633, 287.6472, 287.6313, 287.6155, 287.5996, 287.5835, 287.5676, 
    287.5518, 287.5359, 287.5461, 287.5566, 287.5671, 287.5774, 287.5879, 
    287.5984, 287.6086, 287.6191, 287.6296, 287.6399, 287.6504, 287.6609, 
    287.6689, 287.6748, 287.6807, 287.6865, 287.6924, 287.6982, 287.7041, 
    287.71, 287.7158, 287.7214, 287.7273, 287.7332, 287.739, 287.7344, 
    287.7297, 287.7251, 287.7205, 287.7158, 287.7112, 287.7065, 287.7019, 
    287.6973, 287.6926, 287.688, 287.6833, 287.6794, 287.6763, 287.6731, 
    287.6702, 287.667, 287.6638, 287.6606, 287.6575, 287.6543, 287.6511, 
    287.6479, 287.6448, 287.6416, 287.6387, 287.6355, 287.6326, 287.6296, 
    287.6265, 287.6235, 287.6204, 287.6174, 287.6143, 287.6113, 287.6084, 
    287.6052, 287.5869, 287.5496, 287.5063, 287.4563, 287.397, 287.3262, 
    287.2397, 287.1321, 286.9941, 286.8113, 286.5569, 286.1792, 285.5598, 
    285.3445, 285.1289, 284.9136, 284.6982, 284.4827, 284.2673, 284.0518, 
    283.8364, 283.6208, 283.4055, 283.1899, 282.9746, 282.8506, 282.8179, 
    282.7854, 282.7527, 282.7202, 282.6875, 282.6548, 282.6223, 282.5896, 
    282.5571, 282.5244, 282.4917, 282.4592, 282.4814, 282.5037, 282.5256, 
    282.5479, 282.5701, 282.5923, 282.6145, 282.6367, 282.6587, 282.6809, 
    282.7031, 282.7253, 282.7473, 282.769, 282.7908, 282.8127, 282.8345, 
    282.8562, 282.8779, 282.8997, 282.9216, 282.9434, 282.9651, 282.9868, 
    283.0088, 282.9521, 282.8955, 282.8389, 282.7822, 282.7256, 282.6689, 
    282.6123, 282.5559, 282.4993, 282.4426, 282.386, 282.3293, 282.2615, 
    282.1824, 282.1033, 282.0242, 281.9451, 281.866, 281.7869, 281.7078, 
    281.6287, 281.5496, 281.4705, 281.3914, 281.3123, 281.2544, 281.1965, 
    281.1387, 281.0806, 281.0227, 280.9648, 280.907, 280.8491, 280.7913, 
    280.7332, 280.6753, 280.6174, 280.5503, 280.4739, 280.3977, 280.3213, 
    280.2449, 280.1687, 280.0923, 280.0159, 279.9397, 279.8633, 279.7869, 
    279.7104, 279.6343, 279.6057, 279.5771, 279.5486, 279.52, 279.4917, 
    279.4631, 279.4346, 279.406, 279.3774, 279.3489, 279.3203, 279.292, 
    279.2642, 279.2371, 279.21, 279.1826, 279.1555, 279.1284, 279.1013, 
    279.0742, 279.0471, 279.02, 278.9929, 278.9658, 278.9387,
  284.708, 284.7371, 285.6445, 285.7393, 285.8162, 285.8799, 285.9333, 
    285.979, 286.0186, 286.053, 286.0833, 286.2014, 286.3152, 286.4248, 
    286.5308, 286.6331, 286.7317, 286.8271, 286.9192, 287.0085, 287.095, 
    287.1787, 287.2598, 287.3193, 287.3594, 287.3992, 287.4392, 287.479, 
    287.519, 287.5591, 287.5989, 287.6389, 287.6787, 287.7188, 287.7585, 
    287.7986, 287.7998, 287.801, 287.8022, 287.8035, 287.8047, 287.8059, 
    287.8071, 287.8083, 287.8096, 287.8108, 287.812, 287.8132, 287.8269, 
    287.8528, 287.8787, 287.9043, 287.9302, 287.9561, 287.9819, 288.0078, 
    288.0337, 288.0593, 288.0852, 288.1111, 288.137, 288.1072, 288.0774, 
    288.0476, 288.0178, 287.988, 287.9583, 287.9285, 287.8987, 287.8689, 
    287.8391, 287.8093, 287.7795, 287.7539, 287.7324, 287.7107, 287.6892, 
    287.6675, 287.646, 287.6245, 287.6028, 287.5813, 287.5596, 287.5381, 
    287.5166, 287.4949, 287.5093, 287.5234, 287.5376, 287.5518, 287.5662, 
    287.5803, 287.5945, 287.6086, 287.6228, 287.6372, 287.6514, 287.6655, 
    287.6753, 287.6807, 287.686, 287.6914, 287.6968, 287.7021, 287.7075, 
    287.7129, 287.7183, 287.7236, 287.729, 287.7344, 287.7397, 287.7363, 
    287.7332, 287.7297, 287.7266, 287.7234, 287.72, 287.7168, 287.7136, 
    287.7102, 287.707, 287.7039, 287.7004, 287.6958, 287.6897, 287.6836, 
    287.6775, 287.6714, 287.6653, 287.6592, 287.6531, 287.647, 287.6409, 
    287.6348, 287.6287, 287.6226, 287.626, 287.6294, 287.6326, 287.636, 
    287.6394, 287.6428, 287.6462, 287.6497, 287.6531, 287.6565, 287.6599, 
    287.6631, 287.6511, 287.6204, 287.5852, 287.5442, 287.4956, 287.4375, 
    287.3667, 287.2786, 287.1655, 287.0159, 286.8074, 286.4983, 285.991, 
    285.7539, 285.5168, 285.28, 285.043, 284.8059, 284.5691, 284.332, 
    284.095, 283.8582, 283.6211, 283.384, 283.147, 283.0046, 282.9565, 
    282.9084, 282.8601, 282.812, 282.7639, 282.7158, 282.6677, 282.6196, 
    282.5715, 282.5234, 282.4753, 282.4272, 282.4443, 282.4617, 282.4788, 
    282.4958, 282.5132, 282.5303, 282.5474, 282.5647, 282.5818, 282.5991, 
    282.6162, 282.6333, 282.6509, 282.6687, 282.6865, 282.7043, 282.7222, 
    282.7397, 282.7576, 282.7754, 282.7932, 282.811, 282.8289, 282.8467, 
    282.8645, 282.8113, 282.7578, 282.7046, 282.6514, 282.5981, 282.5447, 
    282.4915, 282.4382, 282.385, 282.3318, 282.2783, 282.2251, 282.1646, 
    282.0964, 282.0283, 281.9604, 281.8923, 281.8245, 281.7563, 281.6882, 
    281.6204, 281.5522, 281.4841, 281.4163, 281.3481, 281.2793, 281.2107, 
    281.1418, 281.0732, 281.0044, 280.9355, 280.8669, 280.7981, 280.7295, 
    280.6606, 280.5918, 280.5232, 280.4524, 280.3794, 280.3066, 280.2336, 
    280.1609, 280.0879, 280.0151, 279.9421, 279.8694, 279.7964, 279.7236, 
    279.6506, 279.5779, 279.5542, 279.5308, 279.5071, 279.4836, 279.46, 
    279.4365, 279.4131, 279.3894, 279.366, 279.3423, 279.3188, 279.2952, 
    279.2676, 279.2358, 279.2041, 279.1724, 279.1406, 279.1089, 279.0771, 
    279.0454, 279.0137, 278.9819, 278.9502, 278.9185, 278.8867,
  284.9302, 284.9563, 285.7854, 285.8633, 285.9255, 285.9766, 286.019, 
    286.0549, 286.0854, 286.1121, 286.1355, 286.252, 286.3667, 286.48, 
    286.5918, 286.7021, 286.811, 286.9185, 287.0247, 287.1294, 287.2329, 
    287.335, 287.436, 287.4993, 287.5256, 287.5522, 287.5786, 287.6052, 
    287.6318, 287.6582, 287.6848, 287.7114, 287.7378, 287.7644, 287.791, 
    287.8174, 287.8184, 287.8193, 287.8203, 287.8213, 287.8223, 287.8232, 
    287.8242, 287.8252, 287.8262, 287.8271, 287.8281, 287.8291, 287.8445, 
    287.8743, 287.9043, 287.9341, 287.9641, 287.9939, 288.0237, 288.0537, 
    288.0835, 288.1135, 288.1433, 288.1731, 288.2031, 288.1704, 288.1377, 
    288.105, 288.0723, 288.0396, 288.0068, 287.9741, 287.9417, 287.9089, 
    287.8762, 287.8435, 287.8108, 287.7808, 287.7537, 287.7263, 287.6992, 
    287.6719, 287.6448, 287.6174, 287.5903, 287.563, 287.5359, 287.5085, 
    287.4814, 287.4541, 287.4722, 287.4902, 287.5081, 287.5261, 287.5442, 
    287.5623, 287.5803, 287.5981, 287.6162, 287.6343, 287.6523, 287.6704, 
    287.6819, 287.6868, 287.6914, 287.6963, 287.7012, 287.7061, 287.7109, 
    287.7158, 287.7207, 287.7256, 287.7305, 287.7354, 287.7402, 287.7383, 
    287.7363, 287.7346, 287.7327, 287.7307, 287.729, 287.7271, 287.7251, 
    287.7231, 287.7214, 287.7195, 287.7175, 287.7122, 287.7031, 287.6941, 
    287.6848, 287.6758, 287.6667, 287.6577, 287.6487, 287.6396, 287.6306, 
    287.6213, 287.6123, 287.6033, 287.613, 287.623, 287.6328, 287.6426, 
    287.6523, 287.6621, 287.6721, 287.6819, 287.6917, 287.7014, 287.7114, 
    287.7212, 287.7153, 287.6914, 287.6638, 287.6318, 287.5942, 287.5488, 
    287.4939, 287.425, 287.3372, 287.2205, 287.0581, 286.8171, 286.4219, 
    286.1633, 285.9048, 285.6462, 285.3877, 285.1292, 284.8708, 284.6123, 
    284.3538, 284.0952, 283.8367, 283.5781, 283.3196, 283.1584, 283.095, 
    283.0312, 282.9678, 282.9041, 282.8406, 282.7769, 282.7134, 282.6497, 
    282.5862, 282.5225, 282.459, 282.3953, 282.4075, 282.4197, 282.4319, 
    282.4441, 282.4561, 282.4683, 282.4805, 282.4927, 282.5049, 282.5171, 
    282.5293, 282.5415, 282.5544, 282.5681, 282.582, 282.5959, 282.6096, 
    282.6235, 282.6372, 282.6511, 282.665, 282.6787, 282.6926, 282.7063, 
    282.7202, 282.6702, 282.6204, 282.5703, 282.5205, 282.4705, 282.4207, 
    282.3706, 282.3208, 282.2708, 282.2207, 282.1709, 282.1208, 282.0674, 
    282.0105, 281.9536, 281.8967, 281.8396, 281.7827, 281.7258, 281.6687, 
    281.6118, 281.5549, 281.4978, 281.4409, 281.384, 281.3044, 281.2249, 
    281.1453, 281.0657, 280.9861, 280.9065, 280.8269, 280.7471, 280.6675, 
    280.5879, 280.5083, 280.4287, 280.3542, 280.2849, 280.2156, 280.146, 
    280.0767, 280.0073, 279.9377, 279.8684, 279.7991, 279.7297, 279.6602, 
    279.5908, 279.5215, 279.5029, 279.4844, 279.4656, 279.447, 279.4285, 
    279.4099, 279.3914, 279.3728, 279.3542, 279.3357, 279.3171, 279.2986, 
    279.2712, 279.2349, 279.1985, 279.1621, 279.1257, 279.0894, 279.053, 
    279.0166, 278.9802, 278.9438, 278.9075, 278.8711, 278.8347,
  285.1086, 285.1382, 285.9636, 286.0195, 286.0647, 286.1018, 286.1331, 
    286.1597, 286.1824, 286.2021, 286.2197, 286.3325, 286.4456, 286.5583, 
    286.6714, 286.7842, 286.8972, 287.0103, 287.123, 287.2361, 287.3489, 
    287.4619, 287.575, 287.6399, 287.6572, 287.6746, 287.6919, 287.7092, 
    287.7266, 287.7439, 287.7612, 287.7786, 287.7959, 287.8132, 287.8306, 
    287.8479, 287.8484, 287.8491, 287.8499, 287.8506, 287.8513, 287.8518, 
    287.8525, 287.8533, 287.854, 287.8545, 287.8552, 287.856, 287.8721, 
    287.9038, 287.9355, 287.9673, 287.999, 288.0305, 288.0623, 288.094, 
    288.1257, 288.1575, 288.1892, 288.2207, 288.2524, 288.2178, 288.1831, 
    288.1484, 288.1135, 288.0789, 288.0442, 288.0095, 287.9749, 287.9399, 
    287.9053, 287.8706, 287.8359, 287.8032, 287.7725, 287.7419, 287.7112, 
    287.6807, 287.6499, 287.6194, 287.5886, 287.5579, 287.5273, 287.4966, 
    287.4661, 287.4353, 287.4561, 287.4768, 287.4973, 287.5181, 287.5388, 
    287.5596, 287.5801, 287.6008, 287.6216, 287.6423, 287.6628, 287.6836, 
    287.6953, 287.698, 287.7007, 287.7034, 287.7063, 287.709, 287.7117, 
    287.7144, 287.717, 287.7197, 287.7224, 287.7251, 287.7278, 287.7275, 
    287.7273, 287.7271, 287.7268, 287.7266, 287.7263, 287.7261, 287.7256, 
    287.7253, 287.7251, 287.7249, 287.7246, 287.719, 287.7083, 287.6973, 
    287.6865, 287.6755, 287.6648, 287.6538, 287.6431, 287.6321, 287.6213, 
    287.6104, 287.5996, 287.5886, 287.6025, 287.6162, 287.6301, 287.6438, 
    287.6577, 287.6714, 287.6853, 287.699, 287.7126, 287.7266, 287.7402, 
    287.7542, 287.7527, 287.7341, 287.7129, 287.688, 287.6587, 287.6235, 
    287.5808, 287.5276, 287.4592, 287.3687, 287.2427, 287.0557, 286.749, 
    286.4753, 286.2017, 285.9277, 285.6541, 285.3804, 285.1067, 284.8328, 
    284.5591, 284.2854, 284.0115, 283.7378, 283.4641, 283.2886, 283.2112, 
    283.134, 283.0566, 282.9795, 282.9021, 282.8247, 282.7476, 282.6702, 
    282.593, 282.5156, 282.4382, 282.3611, 282.3711, 282.3809, 282.3909, 
    282.4009, 282.4109, 282.4207, 282.4307, 282.4407, 282.4507, 282.4607, 
    282.4705, 282.4805, 282.4893, 282.4971, 282.5049, 282.5127, 282.5205, 
    282.5283, 282.5361, 282.5439, 282.5518, 282.5596, 282.5674, 282.5752, 
    282.583, 282.5361, 282.4893, 282.4426, 282.3958, 282.3489, 282.302, 
    282.2554, 282.2085, 282.1616, 282.1147, 282.0681, 282.0212, 281.9744, 
    281.9275, 281.8806, 281.8337, 281.7869, 281.74, 281.6931, 281.6462, 
    281.5994, 281.5525, 281.5056, 281.4587, 281.4119, 281.3237, 281.2358, 
    281.1479, 281.0601, 280.9722, 280.8843, 280.7961, 280.7083, 280.6204, 
    280.5325, 280.4446, 280.3564, 280.2791, 280.2119, 280.1445, 280.0774, 
    280.0103, 279.9431, 279.876, 279.8086, 279.7415, 279.6743, 279.6072, 
    279.54, 279.4729, 279.4565, 279.4404, 279.4243, 279.408, 279.3918, 
    279.3757, 279.3596, 279.3433, 279.3271, 279.311, 279.2949, 279.2786, 
    279.2522, 279.2156, 279.1792, 279.1426, 279.106, 279.0693, 279.0327, 
    278.9961, 278.9595, 278.9231, 278.8865, 278.8499, 278.8132,
  285.1804, 285.2168, 286.2168, 286.2517, 286.2815, 286.3071, 286.3293, 
    286.3486, 286.366, 286.3813, 286.395, 286.4983, 286.6018, 286.7051, 
    286.8086, 286.9119, 287.0154, 287.1187, 287.2222, 287.3254, 287.429, 
    287.5322, 287.6357, 287.696, 287.7134, 287.7305, 287.7478, 287.7651, 
    287.7822, 287.7996, 287.8169, 287.8342, 287.8513, 287.8687, 287.886, 
    287.9031, 287.9036, 287.9038, 287.9041, 287.9045, 287.9048, 287.9053, 
    287.9055, 287.9058, 287.9062, 287.9065, 287.907, 287.9072, 287.9216, 
    287.9504, 287.979, 288.0078, 288.0364, 288.0649, 288.0938, 288.1223, 
    288.1509, 288.1797, 288.2083, 288.2368, 288.2656, 288.2307, 288.196, 
    288.1611, 288.1262, 288.0916, 288.0566, 288.022, 287.9871, 287.9524, 
    287.9175, 287.8828, 287.8479, 287.8159, 287.7866, 287.7573, 287.728, 
    287.6987, 287.6694, 287.6401, 287.6108, 287.5815, 287.5522, 287.5229, 
    287.4937, 287.4646, 287.4854, 287.5063, 287.5273, 287.5481, 287.5691, 
    287.5901, 287.6108, 287.6318, 287.6528, 287.6736, 287.6946, 287.7156, 
    287.7244, 287.7214, 287.7183, 287.7151, 287.7122, 287.709, 287.7061, 
    287.7029, 287.7, 287.6968, 287.6936, 287.6907, 287.6875, 287.6895, 
    287.6912, 287.6931, 287.6948, 287.6968, 287.6987, 287.7004, 287.7024, 
    287.7041, 287.7061, 287.7078, 287.7097, 287.7056, 287.6953, 287.6853, 
    287.675, 287.665, 287.6548, 287.6448, 287.6345, 287.6245, 287.6143, 
    287.6042, 287.594, 287.584, 287.5964, 287.6089, 287.6211, 287.6335, 
    287.646, 287.6584, 287.6709, 287.6831, 287.6956, 287.708, 287.7205, 
    287.7329, 287.7317, 287.7156, 287.6968, 287.6748, 287.6492, 287.6184, 
    287.5808, 287.5339, 287.4741, 287.3945, 287.2839, 287.1199, 286.8506, 
    286.5752, 286.3, 286.0249, 285.7495, 285.4744, 285.199, 284.9238, 
    284.6487, 284.3733, 284.0981, 283.8228, 283.5476, 283.3665, 283.2795, 
    283.1924, 283.1052, 283.0183, 282.9312, 282.8442, 282.7571, 282.6702, 
    282.583, 282.4958, 282.4089, 282.3218, 282.3357, 282.3494, 282.3633, 
    282.377, 282.3909, 282.4045, 282.4182, 282.4321, 282.4458, 282.4597, 
    282.4734, 282.4873, 282.4927, 282.4902, 282.4875, 282.4849, 282.4822, 
    282.4795, 282.4768, 282.4741, 282.4717, 282.469, 282.4663, 282.4636, 
    282.4609, 282.4167, 282.3728, 282.3286, 282.2844, 282.2402, 282.196, 
    282.1519, 282.1079, 282.0637, 282.0195, 281.9753, 281.9312, 281.8896, 
    281.8506, 281.8118, 281.7727, 281.7339, 281.6948, 281.6558, 281.6169, 
    281.5779, 281.5391, 281.5, 281.4609, 281.4221, 281.3313, 281.2405, 
    281.1497, 281.0588, 280.968, 280.8772, 280.7864, 280.6956, 280.6047, 
    280.5139, 280.4233, 280.3325, 280.2532, 280.1855, 280.1179, 280.05, 
    279.9824, 279.9148, 279.8472, 279.7795, 279.7119, 279.644, 279.5764, 
    279.5088, 279.4412, 279.4216, 279.4023, 279.3828, 279.3633, 279.344, 
    279.3245, 279.3052, 279.2856, 279.2664, 279.2468, 279.2275, 279.208, 
    279.1846, 279.1575, 279.1301, 279.103, 279.0757, 279.0486, 279.0212, 
    278.9941, 278.9668, 278.9397, 278.9124, 278.8853, 278.8579,
  285.2732, 285.3174, 286.4136, 286.4417, 286.4663, 286.4885, 286.5083, 
    286.5261, 286.5422, 286.5569, 286.5703, 286.6641, 286.7581, 286.8518, 
    286.9458, 287.0396, 287.1335, 287.2273, 287.3213, 287.415, 287.509, 
    287.6028, 287.6965, 287.7522, 287.7693, 287.7866, 287.8037, 287.8208, 
    287.8381, 287.8552, 287.8726, 287.8896, 287.907, 287.9241, 287.9412, 
    287.9585, 287.9585, 287.9585, 287.9585, 287.9585, 287.9585, 287.9585, 
    287.9585, 287.9585, 287.9585, 287.9585, 287.9585, 287.9585, 287.9714, 
    287.9971, 288.0225, 288.0481, 288.0737, 288.0994, 288.125, 288.1506, 
    288.1763, 288.2019, 288.2273, 288.2529, 288.2786, 288.2437, 288.2087, 
    288.1738, 288.1392, 288.1042, 288.0693, 288.0344, 287.9995, 287.9646, 
    287.9297, 287.8948, 287.8599, 287.8286, 287.8005, 287.7727, 287.7449, 
    287.7168, 287.689, 287.6611, 287.6333, 287.6052, 287.5774, 287.5496, 
    287.5215, 287.4937, 287.5149, 287.5359, 287.5571, 287.5781, 287.5994, 
    287.6206, 287.6416, 287.6628, 287.6838, 287.7051, 287.7263, 287.7473, 
    287.7534, 287.7446, 287.7358, 287.7271, 287.718, 287.7092, 287.7004, 
    287.6917, 287.6826, 287.6738, 287.665, 287.6562, 287.6472, 287.6511, 
    287.6553, 287.6592, 287.6631, 287.667, 287.6709, 287.675, 287.679, 
    287.6829, 287.6868, 287.6907, 287.6948, 287.6919, 287.6826, 287.6731, 
    287.6638, 287.6543, 287.645, 287.6355, 287.6262, 287.6169, 287.6074, 
    287.5981, 287.5886, 287.5793, 287.5903, 287.6013, 287.6123, 287.6233, 
    287.6343, 287.6455, 287.6565, 287.6675, 287.6785, 287.6895, 287.7004, 
    287.7117, 287.7107, 287.6968, 287.6807, 287.6619, 287.6396, 287.6133, 
    287.5808, 287.5405, 287.4888, 287.4204, 287.3252, 287.1838, 286.9519, 
    286.6753, 286.3984, 286.1218, 285.845, 285.5684, 285.2915, 285.0149, 
    284.738, 284.4614, 284.1846, 283.908, 283.6311, 283.4443, 283.3477, 
    283.2507, 283.1541, 283.0571, 282.9604, 282.8635, 282.7668, 282.6699, 
    282.573, 282.4763, 282.3794, 282.2827, 282.3003, 282.3179, 282.3354, 
    282.353, 282.3706, 282.3882, 282.406, 282.4236, 282.4412, 282.4587, 
    282.4763, 282.4939, 282.4961, 282.4832, 282.47, 282.4568, 282.4438, 
    282.4307, 282.4175, 282.4045, 282.3914, 282.3784, 282.3652, 282.3521, 
    282.3391, 282.2976, 282.2561, 282.2146, 282.1731, 282.1316, 282.0901, 
    282.0486, 282.0071, 281.9656, 281.9243, 281.8828, 281.8413, 281.8049, 
    281.7739, 281.7429, 281.7119, 281.6807, 281.6497, 281.6187, 281.5876, 
    281.5566, 281.5254, 281.4944, 281.4634, 281.4324, 281.3386, 281.2451, 
    281.1514, 281.0576, 280.9641, 280.8704, 280.7766, 280.6829, 280.5894, 
    280.4956, 280.4019, 280.3083, 280.2273, 280.1592, 280.0911, 280.0229, 
    279.9548, 279.8865, 279.8184, 279.7502, 279.6821, 279.614, 279.5457, 
    279.4775, 279.4094, 279.3867, 279.364, 279.3413, 279.3188, 279.2961, 
    279.2734, 279.2507, 279.228, 279.2053, 279.1826, 279.1602, 279.1375, 
    279.1172, 279.0994, 279.0813, 279.0635, 279.0457, 279.0278, 279.01, 
    278.9919, 278.9741, 278.9563, 278.9385, 278.9207, 278.9028,
  285.397, 285.4504, 286.5713, 286.5999, 286.626, 286.6499, 286.6721, 
    286.6926, 286.7117, 286.7292, 286.7456, 286.8301, 286.9143, 286.9985, 
    287.083, 287.1672, 287.2517, 287.3359, 287.4202, 287.5046, 287.5889, 
    287.6731, 287.7576, 287.8083, 287.8254, 287.8425, 287.8596, 287.8767, 
    287.8938, 287.9109, 287.9282, 287.9453, 287.9624, 287.9795, 287.9966, 
    288.0137, 288.0134, 288.0132, 288.0127, 288.0125, 288.0122, 288.0117, 
    288.0115, 288.0112, 288.0107, 288.0105, 288.0103, 288.0098, 288.021, 
    288.0435, 288.0662, 288.0886, 288.1111, 288.1338, 288.1562, 288.179, 
    288.2014, 288.2239, 288.2466, 288.269, 288.2917, 288.2566, 288.2217, 
    288.1868, 288.1519, 288.1167, 288.0818, 288.0469, 288.0117, 287.9768, 
    287.9419, 287.907, 287.8718, 287.8411, 287.8147, 287.7881, 287.7615, 
    287.7351, 287.7085, 287.6819, 287.6555, 287.6289, 287.6023, 287.5759, 
    287.5493, 287.5229, 287.5442, 287.5657, 287.5869, 287.6084, 287.6296, 
    287.6511, 287.6724, 287.6938, 287.7151, 287.7366, 287.7578, 287.7793, 
    287.7825, 287.7678, 287.7532, 287.7388, 287.7241, 287.7095, 287.6948, 
    287.6802, 287.6655, 287.6509, 287.6362, 287.6216, 287.6069, 287.613, 
    287.6191, 287.6252, 287.6313, 287.6372, 287.6433, 287.6494, 287.6555, 
    287.6616, 287.6677, 287.6736, 287.6797, 287.6785, 287.6697, 287.6611, 
    287.6526, 287.6438, 287.6353, 287.6265, 287.6179, 287.6091, 287.6006, 
    287.5918, 287.5833, 287.5745, 287.5842, 287.5938, 287.6035, 287.613, 
    287.6228, 287.6323, 287.6421, 287.6516, 287.6614, 287.6709, 287.6807, 
    287.6904, 287.6899, 287.6782, 287.6646, 287.6489, 287.6301, 287.6079, 
    287.5808, 287.5471, 287.5037, 287.4463, 287.3665, 287.2478, 287.0535, 
    286.7751, 286.4968, 286.2188, 285.9404, 285.6624, 285.384, 285.106, 
    284.8276, 284.5493, 284.2712, 283.9929, 283.7148, 283.5225, 283.4158, 
    283.3093, 283.2026, 283.0959, 282.9895, 282.8828, 282.7764, 282.6697, 
    282.5632, 282.4565, 282.3501, 282.2434, 282.2649, 282.2864, 282.3079, 
    282.3291, 282.3506, 282.3721, 282.3936, 282.4148, 282.4363, 282.4578, 
    282.4792, 282.5005, 282.4995, 282.4761, 282.4524, 282.429, 282.4053, 
    282.3818, 282.3584, 282.3347, 282.3113, 282.2876, 282.2642, 282.2405, 
    282.217, 282.1782, 282.1394, 282.1006, 282.0618, 282.0229, 281.9841, 
    281.9453, 281.9065, 281.8677, 281.8289, 281.79, 281.7512, 281.7202, 
    281.6973, 281.6741, 281.6509, 281.6277, 281.6045, 281.5815, 281.5583, 
    281.5352, 281.512, 281.489, 281.4658, 281.4426, 281.3462, 281.2495, 
    281.1531, 281.0564, 280.96, 280.8633, 280.7668, 280.6704, 280.5737, 
    280.4773, 280.3806, 280.2842, 280.2017, 280.1328, 280.0642, 279.9956, 
    279.927, 279.8584, 279.7896, 279.7209, 279.6523, 279.5837, 279.5151, 
    279.4463, 279.3777, 279.3518, 279.3259, 279.3, 279.2742, 279.248, 
    279.2222, 279.1963, 279.1704, 279.1445, 279.1187, 279.0928, 279.0667, 
    279.0496, 279.041, 279.0325, 279.0239, 279.0156, 279.0071, 278.9985, 
    278.99, 278.9814, 278.9729, 278.9646, 278.9561, 278.9475,
  285.5715, 285.6355, 286.7002, 286.7336, 286.7651, 286.7947, 286.8228, 
    286.8494, 286.8745, 286.8984, 286.9209, 286.9958, 287.0706, 287.1453, 
    287.2202, 287.2949, 287.3696, 287.4446, 287.5193, 287.594, 287.6689, 
    287.7437, 287.8184, 287.8643, 287.8813, 287.8984, 287.9155, 287.9326, 
    287.9497, 287.9668, 287.9836, 288.0007, 288.0178, 288.0349, 288.052, 
    288.0691, 288.0684, 288.0676, 288.0671, 288.0664, 288.0657, 288.0652, 
    288.0645, 288.0637, 288.0632, 288.0625, 288.0618, 288.061, 288.0706, 
    288.0901, 288.1096, 288.1292, 288.1487, 288.1682, 288.1877, 288.2073, 
    288.2266, 288.2461, 288.2656, 288.2852, 288.3047, 288.2698, 288.2346, 
    288.1995, 288.1646, 288.1294, 288.0942, 288.0593, 288.0242, 287.989, 
    287.9541, 287.9189, 287.8838, 287.8538, 287.8286, 287.8035, 287.7783, 
    287.7532, 287.728, 287.7029, 287.6777, 287.6526, 287.6274, 287.6023, 
    287.5771, 287.552, 287.5735, 287.5952, 287.6167, 287.6384, 287.6599, 
    287.6816, 287.7031, 287.7246, 287.7463, 287.7678, 287.7896, 287.811, 
    287.8115, 287.7913, 287.7708, 287.7505, 287.73, 287.7095, 287.6892, 
    287.6687, 287.6484, 287.6279, 287.6074, 287.5872, 287.5667, 287.575, 
    287.583, 287.5913, 287.5994, 287.6077, 287.6157, 287.624, 287.6321, 
    287.6404, 287.6484, 287.6567, 287.6648, 287.665, 287.657, 287.6492, 
    287.6411, 287.6333, 287.6252, 287.6174, 287.6094, 287.6016, 287.5935, 
    287.5857, 287.5776, 287.5698, 287.5781, 287.5864, 287.5947, 287.6028, 
    287.6111, 287.6194, 287.6277, 287.636, 287.6443, 287.6526, 287.6609, 
    287.6689, 287.6689, 287.6594, 287.6484, 287.6357, 287.6208, 287.6028, 
    287.5808, 287.5535, 287.5186, 287.4722, 287.4077, 287.3118, 287.1548, 
    286.875, 286.5955, 286.3157, 286.0359, 285.7563, 285.4766, 285.1968, 
    284.9172, 284.6375, 284.3577, 284.0781, 283.7983, 283.6003, 283.4839, 
    283.3677, 283.2512, 283.135, 283.0186, 282.9023, 282.7859, 282.6697, 
    282.5532, 282.437, 282.3206, 282.2043, 282.2295, 282.2549, 282.28, 
    282.3054, 282.3306, 282.3557, 282.3811, 282.4062, 282.4316, 282.4568, 
    282.4819, 282.5073, 282.5029, 282.469, 282.4351, 282.4009, 282.3669, 
    282.333, 282.2991, 282.2649, 282.231, 282.197, 282.1631, 282.1289, 
    282.095, 282.0588, 282.0227, 281.9866, 281.9504, 281.9143, 281.8782, 
    281.842, 281.8059, 281.7698, 281.7336, 281.6975, 281.6614, 281.6355, 
    281.6204, 281.6052, 281.5898, 281.5747, 281.5596, 281.5442, 281.5291, 
    281.5139, 281.4985, 281.4834, 281.468, 281.4529, 281.3535, 281.2542, 
    281.1548, 281.0552, 280.9558, 280.8564, 280.7571, 280.6577, 280.5583, 
    280.4587, 280.3594, 280.26, 280.1758, 280.1067, 280.0376, 279.9683, 
    279.8992, 279.8301, 279.761, 279.6917, 279.6226, 279.5535, 279.4844, 
    279.4153, 279.3459, 279.3169, 279.2878, 279.2585, 279.2295, 279.2002, 
    279.1711, 279.1418, 279.1128, 279.0835, 279.0544, 279.0254, 278.9961, 
    278.9819, 278.9829, 278.9836, 278.9846, 278.9854, 278.9863, 278.9871, 
    278.988, 278.9888, 278.9897, 278.9905, 278.9915, 278.9922,
  286.7222, 286.7659, 286.8079, 286.8481, 286.8875, 286.925, 286.9617, 
    286.9971, 287.0312, 287.0642, 287.0964, 287.1616, 287.2268, 287.292, 
    287.3574, 287.4226, 287.4878, 287.553, 287.6184, 287.6836, 287.7488, 
    287.8142, 287.8794, 287.9204, 287.9375, 287.9543, 287.9714, 287.9885, 
    288.0054, 288.0225, 288.0393, 288.0564, 288.0732, 288.0903, 288.1074, 
    288.1243, 288.1233, 288.1223, 288.1213, 288.1204, 288.1194, 288.1184, 
    288.1174, 288.1165, 288.1155, 288.1145, 288.1135, 288.1125, 288.1201, 
    288.1367, 288.1531, 288.1697, 288.186, 288.2026, 288.219, 288.2354, 
    288.252, 288.2683, 288.2849, 288.3013, 288.3179, 288.2827, 288.2476, 
    288.2124, 288.1772, 288.1421, 288.1069, 288.0718, 288.0366, 288.0015, 
    287.9663, 287.9312, 287.896, 287.8665, 287.8425, 287.8188, 287.7952, 
    287.7712, 287.7476, 287.7239, 287.7, 287.6763, 287.6526, 287.6287, 
    287.605, 287.5813, 287.603, 287.6248, 287.6467, 287.6685, 287.6902, 
    287.7122, 287.7339, 287.7556, 287.7773, 287.7993, 287.821, 287.8428, 
    287.8406, 287.8145, 287.7883, 287.7622, 287.7358, 287.7097, 287.6836, 
    287.6575, 287.6311, 287.605, 287.5789, 287.5525, 287.5264, 287.5366, 
    287.5469, 287.5574, 287.5676, 287.5779, 287.5881, 287.5984, 287.6086, 
    287.6189, 287.6294, 287.6396, 287.6499, 287.6514, 287.6443, 287.637, 
    287.6299, 287.6226, 287.6155, 287.6082, 287.6011, 287.5938, 287.5867, 
    287.5793, 287.5723, 287.5652, 287.572, 287.5789, 287.5857, 287.5925, 
    287.5996, 287.6064, 287.6133, 287.6201, 287.6272, 287.634, 287.6409, 
    287.6477, 287.6479, 287.6406, 287.6323, 287.6228, 287.6113, 287.5977, 
    287.5808, 287.5601, 287.5334, 287.498, 287.449, 287.376, 287.2561, 
    286.9751, 286.6938, 286.4126, 286.1313, 285.8503, 285.5691, 285.2878, 
    285.0066, 284.7253, 284.4443, 284.1631, 283.8818, 283.6782, 283.552, 
    283.426, 283.3, 283.1738, 283.0479, 282.9216, 282.7957, 282.6694, 
    282.5435, 282.4172, 282.2913, 282.165, 282.1941, 282.2234, 282.2524, 
    282.2815, 282.3105, 282.3396, 282.3687, 282.3977, 282.4268, 282.4558, 
    282.4849, 282.5139, 282.5063, 282.4619, 282.4175, 282.373, 282.3286, 
    282.2842, 282.2397, 282.1953, 282.1509, 282.1064, 282.062, 282.0176, 
    281.9731, 281.9395, 281.906, 281.8726, 281.8391, 281.8057, 281.7722, 
    281.7388, 281.7053, 281.6716, 281.6382, 281.6047, 281.5713, 281.551, 
    281.5437, 281.5364, 281.5291, 281.5217, 281.5144, 281.5071, 281.4998, 
    281.4924, 281.4851, 281.4778, 281.4705, 281.4631, 281.3608, 281.2585, 
    281.1562, 281.0542, 280.9519, 280.8496, 280.7473, 280.645, 280.5427, 
    280.4404, 280.3381, 280.2358, 280.1499, 280.0803, 280.0107, 279.9412, 
    279.8713, 279.8018, 279.7322, 279.6626, 279.593, 279.5232, 279.4536, 
    279.384, 279.3145, 279.282, 279.2495, 279.217, 279.1848, 279.1523, 
    279.1199, 279.0876, 279.0552, 279.0227, 278.9902, 278.958, 278.9255, 
    278.9143, 278.9246, 278.9348, 278.9451, 278.9553, 278.9656, 278.9756, 
    278.9858, 278.9961, 279.0063, 279.0166, 279.0269, 279.0369,
  286.7991, 286.8491, 286.8987, 286.9475, 286.9958, 287.0432, 287.0901, 
    287.1365, 287.1821, 287.2273, 287.2717, 287.3274, 287.3831, 287.439, 
    287.4946, 287.5503, 287.606, 287.6616, 287.7173, 287.7732, 287.8289, 
    287.8845, 287.9402, 287.9766, 287.9934, 288.0105, 288.0273, 288.0442, 
    288.0613, 288.0781, 288.095, 288.1121, 288.1289, 288.1458, 288.1626, 
    288.1797, 288.1782, 288.177, 288.1755, 288.1743, 288.1731, 288.1716, 
    288.1704, 288.1689, 288.1677, 288.1665, 288.165, 288.1638, 288.1697, 
    288.1831, 288.1965, 288.21, 288.2234, 288.2368, 288.2502, 288.2637, 
    288.2771, 288.2905, 288.304, 288.3174, 288.3308, 288.2957, 288.2603, 
    288.2251, 288.1899, 288.1545, 288.1194, 288.0842, 288.0488, 288.0137, 
    287.9783, 287.9431, 287.908, 287.8792, 287.8567, 287.8342, 287.8118, 
    287.7896, 287.7671, 287.7446, 287.7224, 287.7, 287.6775, 287.6553, 
    287.6328, 287.6104, 287.6323, 287.6545, 287.6765, 287.6985, 287.7205, 
    287.7424, 287.7646, 287.7866, 287.8086, 287.8306, 287.8528, 287.8748, 
    287.8699, 287.8379, 287.8059, 287.7739, 287.7419, 287.71, 287.678, 
    287.646, 287.614, 287.582, 287.55, 287.5181, 287.4861, 287.4985, 287.511, 
    287.5232, 287.5356, 287.5481, 287.5605, 287.573, 287.5852, 287.5977, 
    287.6101, 287.6226, 287.635, 287.6379, 287.6313, 287.625, 287.6184, 
    287.6121, 287.6055, 287.5991, 287.5928, 287.5862, 287.5798, 287.5732, 
    287.5669, 287.5603, 287.5659, 287.5713, 287.5769, 287.5825, 287.5879, 
    287.5935, 287.5989, 287.6045, 287.6099, 287.6155, 287.6211, 287.6265, 
    287.627, 287.6221, 287.6165, 287.6096, 287.6018, 287.5923, 287.5808, 
    287.5667, 287.5483, 287.5239, 287.4902, 287.4399, 287.3577, 287.075, 
    286.7922, 286.5095, 286.2268, 285.9443, 285.6616, 285.3789, 285.0962, 
    284.8135, 284.5308, 284.248, 283.9653, 283.7561, 283.6204, 283.4844, 
    283.3486, 283.2126, 283.0769, 282.9412, 282.8052, 282.6694, 282.5334, 
    282.3977, 282.2617, 282.126, 282.1589, 282.1917, 282.2246, 282.2576, 
    282.2905, 282.3232, 282.3562, 282.3892, 282.4221, 282.4548, 282.4878, 
    282.5208, 282.5098, 282.4548, 282.3999, 282.345, 282.29, 282.2354, 
    282.1804, 282.1255, 282.0706, 282.0156, 281.9609, 281.906, 281.8511, 
    281.8203, 281.7896, 281.7585, 281.7278, 281.697, 281.6663, 281.6355, 
    281.6045, 281.5737, 281.543, 281.5122, 281.4814, 281.4663, 281.4668, 
    281.4675, 281.468, 281.4688, 281.4692, 281.47, 281.4705, 281.4709, 
    281.4717, 281.4722, 281.4729, 281.4734, 281.3684, 281.2632, 281.158, 
    281.053, 280.9478, 280.8425, 280.7375, 280.6323, 280.5271, 280.4221, 
    280.3169, 280.2117, 280.124, 280.054, 279.9839, 279.9138, 279.8438, 
    279.7734, 279.7034, 279.6333, 279.5632, 279.4932, 279.4229, 279.3528, 
    279.2827, 279.2471, 279.2114, 279.1758, 279.1401, 279.1045, 279.0688, 
    279.0332, 278.9976, 278.9619, 278.9263, 278.8906, 278.855, 278.8469, 
    278.8665, 278.886, 278.9055, 278.925, 278.9446, 278.9644, 278.9839, 
    279.0034, 279.0229, 279.0425, 279.062, 279.0818,
  286.8643, 286.9192, 286.9739, 287.0288, 287.0837, 287.1384, 287.1934, 
    287.248, 287.303, 287.3577, 287.4126, 287.4609, 287.5095, 287.5581, 
    287.6064, 287.655, 287.7034, 287.752, 287.8003, 287.8489, 287.8972, 
    287.9458, 287.9941, 288.0269, 288.0437, 288.0605, 288.0771, 288.094, 
    288.1108, 288.1274, 288.1443, 288.1611, 288.1777, 288.1946, 288.2114, 
    288.2283, 288.2256, 288.2229, 288.22, 288.2173, 288.2146, 288.2119, 
    288.2092, 288.2065, 288.2039, 288.2012, 288.1985, 288.1958, 288.2004, 
    288.2122, 288.2241, 288.2358, 288.2476, 288.2595, 288.2712, 288.283, 
    288.2949, 288.3066, 288.3186, 288.3303, 288.342, 288.3076, 288.2732, 
    288.2388, 288.2043, 288.1699, 288.1355, 288.1011, 288.0667, 288.0322, 
    287.9978, 287.9634, 287.929, 287.9004, 287.8774, 287.8545, 287.8318, 
    287.8088, 287.7861, 287.7632, 287.7402, 287.7175, 287.6946, 287.6716, 
    287.6489, 287.626, 287.647, 287.668, 287.689, 287.71, 287.731, 287.752, 
    287.7729, 287.7939, 287.8149, 287.8359, 287.8569, 287.8779, 287.8708, 
    287.8362, 287.8013, 287.7664, 287.7314, 287.6968, 287.6619, 287.627, 
    287.592, 287.5574, 287.5225, 287.4875, 287.4526, 287.467, 287.4814, 
    287.4956, 287.51, 287.5244, 287.5386, 287.553, 287.5674, 287.5815, 
    287.5959, 287.6104, 287.6245, 287.6287, 287.6223, 287.616, 287.6096, 
    287.6033, 287.5969, 287.5906, 287.5842, 287.5779, 287.5715, 287.5654, 
    287.5591, 287.5527, 287.5569, 287.561, 287.5654, 287.5696, 287.5737, 
    287.5781, 287.5823, 287.5864, 287.5908, 287.595, 287.5991, 287.6033, 
    287.6045, 287.6023, 287.5999, 287.5969, 287.5938, 287.5896, 287.585, 
    287.5789, 287.5715, 287.562, 287.5491, 287.5308, 287.4336, 287.1484, 
    286.865, 286.583, 286.3025, 286.0237, 285.7461, 285.47, 285.1956, 
    284.9224, 284.6506, 284.3804, 284.1116, 283.9043, 283.7576, 283.6106, 
    283.4639, 283.3171, 283.1702, 283.0234, 282.8767, 282.7297, 282.583, 
    282.4363, 282.2896, 282.1426, 282.1738, 282.2048, 282.2358, 282.2668, 
    282.2981, 282.3291, 282.3601, 282.3914, 282.4224, 282.4534, 282.4846, 
    282.5156, 282.4995, 282.4363, 282.3733, 282.3101, 282.2468, 282.1836, 
    282.1204, 282.0574, 281.9941, 281.9309, 281.8677, 281.8047, 281.7415, 
    281.7146, 281.688, 281.6611, 281.6345, 281.6077, 281.5811, 281.5542, 
    281.5276, 281.5007, 281.4739, 281.4473, 281.4204, 281.4089, 281.4126, 
    281.4163, 281.4197, 281.4233, 281.427, 281.4307, 281.4341, 281.4377, 
    281.4414, 281.4451, 281.4487, 281.4521, 281.3472, 281.2419, 281.1367, 
    281.0317, 280.9265, 280.8213, 280.7163, 280.6111, 280.5059, 280.4009, 
    280.2957, 280.1904, 280.1047, 280.0386, 279.9722, 279.906, 279.8396, 
    279.7734, 279.707, 279.6409, 279.5745, 279.5083, 279.4419, 279.3757, 
    279.3093, 279.2659, 279.2224, 279.1787, 279.1353, 279.0918, 279.0481, 
    279.0046, 278.9612, 278.9177, 278.874, 278.8306, 278.7871, 278.7788, 
    278.8057, 278.8325, 278.8594, 278.8862, 278.9131, 278.9399, 278.9668, 
    278.9937, 279.0208, 279.0476, 279.0745, 279.1013,
  286.9309, 286.9846, 287.0383, 287.092, 287.1455, 287.1992, 287.2529, 
    287.3066, 287.3604, 287.4138, 287.4675, 287.5146, 287.5615, 287.6084, 
    287.6555, 287.7024, 287.7493, 287.7964, 287.8433, 287.8901, 287.9373, 
    287.9841, 288.0312, 288.0627, 288.0793, 288.0957, 288.1121, 288.1284, 
    288.145, 288.1614, 288.1777, 288.1941, 288.2107, 288.2271, 288.2434, 
    288.2598, 288.2532, 288.2466, 288.24, 288.2334, 288.2268, 288.22, 
    288.2134, 288.2068, 288.2002, 288.1936, 288.187, 288.1804, 288.1838, 
    288.1978, 288.2114, 288.2251, 288.2388, 288.2527, 288.2664, 288.28, 
    288.2937, 288.3076, 288.3213, 288.335, 288.3489, 288.3174, 288.2861, 
    288.2546, 288.2234, 288.1921, 288.1606, 288.1294, 288.0981, 288.0667, 
    288.0354, 288.0042, 287.9727, 287.9431, 287.915, 287.8872, 287.8594, 
    287.8313, 287.8035, 287.7756, 287.7476, 287.7197, 287.6917, 287.6638, 
    287.636, 287.6079, 287.6248, 287.6416, 287.6584, 287.6753, 287.6919, 
    287.7087, 287.7256, 287.7424, 287.7593, 287.7761, 287.793, 287.8096, 
    287.8027, 287.7722, 287.7417, 287.7112, 287.6807, 287.6501, 287.6196, 
    287.5891, 287.5586, 287.5281, 287.4976, 287.467, 287.4365, 287.4524, 
    287.4683, 287.4839, 287.4998, 287.5154, 287.5312, 287.5469, 287.5627, 
    287.5786, 287.5942, 287.6101, 287.6257, 287.6299, 287.6221, 287.6145, 
    287.6067, 287.5991, 287.5916, 287.5837, 287.5762, 287.5684, 287.5608, 
    287.553, 287.5454, 287.5376, 287.5408, 287.5439, 287.5471, 287.5503, 
    287.5535, 287.5566, 287.5598, 287.563, 287.5662, 287.5693, 287.5725, 
    287.5757, 287.5781, 287.5803, 287.583, 287.5857, 287.5891, 287.5928, 
    287.5969, 287.6021, 287.6079, 287.6152, 287.624, 287.6353, 287.4478, 
    287.1575, 286.875, 286.5999, 286.3318, 286.0708, 285.8162, 285.5681, 
    285.3262, 285.0901, 284.8599, 284.635, 284.4153, 284.2271, 284.0664, 
    283.9058, 283.7451, 283.5842, 283.4236, 283.2629, 283.1021, 282.9414, 
    282.7808, 282.6199, 282.4592, 282.2986, 282.3137, 282.3289, 282.3442, 
    282.3594, 282.3745, 282.3899, 282.405, 282.4202, 282.4353, 282.4507, 
    282.4658, 282.481, 282.4556, 282.3894, 282.3235, 282.2573, 282.1912, 
    282.125, 282.0591, 281.9929, 281.9268, 281.8608, 281.7947, 281.7285, 
    281.6626, 281.6433, 281.624, 281.605, 281.5857, 281.5667, 281.5474, 
    281.5283, 281.509, 281.4897, 281.4707, 281.4514, 281.4324, 281.4199, 
    281.4143, 281.4087, 281.4031, 281.3975, 281.3918, 281.3862, 281.3806, 
    281.375, 281.3694, 281.3638, 281.3582, 281.3525, 281.2544, 281.1565, 
    281.0583, 280.9604, 280.8625, 280.7644, 280.6665, 280.5684, 280.4705, 
    280.3723, 280.2744, 280.1763, 280.1016, 280.0498, 279.9983, 279.9465, 
    279.8948, 279.8433, 279.7915, 279.7397, 279.688, 279.6365, 279.5847, 
    279.533, 279.4814, 279.4185, 279.3555, 279.2925, 279.2297, 279.1667, 
    279.1038, 279.0408, 278.9778, 278.915, 278.8521, 278.7891, 278.7261, 
    278.7092, 278.7383, 278.7673, 278.7964, 278.8254, 278.8547, 278.8838, 
    278.9128, 278.9419, 278.9709, 279, 279.0291, 279.0581,
  286.9976, 287.05, 287.1025, 287.155, 287.2075, 287.26, 287.3125, 287.365, 
    287.4175, 287.4702, 287.5227, 287.5681, 287.6135, 287.6589, 287.7043, 
    287.7498, 287.7954, 287.8408, 287.8862, 287.9316, 287.9771, 288.0225, 
    288.0681, 288.0989, 288.1147, 288.1309, 288.147, 288.1631, 288.1792, 
    288.1951, 288.2112, 288.2273, 288.2434, 288.2593, 288.2754, 288.2915, 
    288.281, 288.2705, 288.2598, 288.2493, 288.2388, 288.2283, 288.2175, 
    288.207, 288.1965, 288.186, 288.1753, 288.1648, 288.1675, 288.1831, 
    288.1987, 288.2144, 288.23, 288.2456, 288.2615, 288.2771, 288.2927, 
    288.3083, 288.324, 288.3398, 288.3555, 288.3271, 288.2988, 288.2708, 
    288.2424, 288.2141, 288.186, 288.1577, 288.1294, 288.1013, 288.073, 
    288.0447, 288.0164, 287.9858, 287.9529, 287.9199, 287.887, 287.8538, 
    287.8208, 287.7878, 287.7549, 287.7219, 287.689, 287.656, 287.6228, 
    287.5898, 287.6025, 287.6152, 287.6277, 287.6404, 287.6531, 287.6658, 
    287.6782, 287.6909, 287.7036, 287.7163, 287.7288, 287.7415, 287.7346, 
    287.7085, 287.6824, 287.6562, 287.6299, 287.6038, 287.5776, 287.5515, 
    287.5251, 287.499, 287.4729, 287.4468, 287.4204, 287.4377, 287.4548, 
    287.4722, 287.4893, 287.5066, 287.5237, 287.541, 287.5581, 287.5754, 
    287.5925, 287.6099, 287.627, 287.6311, 287.6221, 287.613, 287.604, 
    287.595, 287.5859, 287.5769, 287.5679, 287.5588, 287.5498, 287.5408, 
    287.5317, 287.5227, 287.5247, 287.5269, 287.5291, 287.531, 287.5332, 
    287.5352, 287.5374, 287.5393, 287.5415, 287.5435, 287.5457, 287.5479, 
    287.552, 287.5591, 287.5669, 287.5754, 287.585, 287.5955, 287.6072, 
    287.6204, 287.6355, 287.6528, 287.6729, 287.6963, 287.4666, 287.1689, 
    286.8872, 286.6201, 286.3665, 286.1255, 285.896, 285.6772, 285.4688, 
    285.2695, 285.0789, 284.8965, 284.7219, 284.55, 284.3755, 284.2007, 
    284.0261, 283.8516, 283.6768, 283.5022, 283.3276, 283.1531, 282.9783, 
    282.8037, 282.6292, 282.4543, 282.4539, 282.4531, 282.4524, 282.4517, 
    282.4512, 282.4504, 282.4497, 282.4492, 282.4485, 282.4478, 282.447, 
    282.4465, 282.4116, 282.3425, 282.2737, 282.2046, 282.1355, 282.0667, 
    281.9976, 281.9285, 281.8596, 281.7905, 281.7217, 281.6526, 281.5835, 
    281.572, 281.5603, 281.5486, 281.5371, 281.5254, 281.5139, 281.5022, 
    281.4905, 281.479, 281.4673, 281.4558, 281.4441, 281.4309, 281.416, 
    281.4011, 281.3862, 281.3713, 281.3567, 281.3418, 281.3269, 281.312, 
    281.2971, 281.2825, 281.2676, 281.2527, 281.1619, 281.071, 280.98, 
    280.8892, 280.7983, 280.7075, 280.6167, 280.5256, 280.4348, 280.344, 
    280.2532, 280.1624, 280.0984, 280.0613, 280.0242, 279.9871, 279.95, 
    279.9128, 279.8757, 279.8389, 279.8018, 279.7646, 279.7275, 279.6904, 
    279.6533, 279.571, 279.4888, 279.4065, 279.324, 279.2417, 279.1594, 
    279.0769, 278.9946, 278.9124, 278.8301, 278.7476, 278.6653, 278.6396, 
    278.6711, 278.7024, 278.7336, 278.7649, 278.7961, 278.8274, 278.8586, 
    278.8899, 278.9214, 278.9526, 278.9839, 279.0151,
  287.064, 287.1155, 287.1667, 287.2183, 287.2695, 287.3208, 287.3723, 
    287.4236, 287.4749, 287.5264, 287.5776, 287.6216, 287.6655, 287.7095, 
    287.7534, 287.7974, 287.8413, 287.8853, 287.9292, 287.9731, 288.0171, 
    288.061, 288.105, 288.1348, 288.1504, 288.1663, 288.1819, 288.1975, 
    288.2134, 288.229, 288.2446, 288.2603, 288.2761, 288.2917, 288.3074, 
    288.3232, 288.3086, 288.2942, 288.2798, 288.2651, 288.2507, 288.2363, 
    288.2217, 288.2073, 288.1926, 288.1782, 288.1638, 288.1492, 288.1509, 
    288.1685, 288.186, 288.2036, 288.2212, 288.2388, 288.2563, 288.2742, 
    288.2917, 288.3093, 288.3269, 288.3445, 288.3621, 288.3369, 288.3118, 
    288.2866, 288.2615, 288.2363, 288.2112, 288.186, 288.1609, 288.1357, 
    288.1106, 288.0854, 288.0603, 288.0286, 287.9905, 287.9524, 287.9143, 
    287.8765, 287.8384, 287.8003, 287.7622, 287.7241, 287.686, 287.6479, 
    287.6099, 287.5718, 287.5803, 287.5886, 287.5972, 287.6057, 287.614, 
    287.6226, 287.6311, 287.6394, 287.6479, 287.6562, 287.6648, 287.6733, 
    287.6665, 287.6448, 287.6228, 287.6011, 287.5791, 287.5574, 287.5354, 
    287.5137, 287.4917, 287.47, 287.448, 287.4263, 287.4043, 287.4231, 
    287.4417, 287.4604, 287.479, 287.4976, 287.5164, 287.5349, 287.5537, 
    287.5723, 287.5911, 287.6096, 287.6282, 287.6323, 287.6221, 287.6116, 
    287.6013, 287.5908, 287.5803, 287.5701, 287.5596, 287.5493, 287.5388, 
    287.5286, 287.5181, 287.5076, 287.5088, 287.5098, 287.5107, 287.5117, 
    287.5127, 287.5139, 287.5149, 287.5159, 287.5168, 287.5178, 287.519, 
    287.52, 287.5264, 287.5386, 287.5518, 287.5659, 287.5811, 287.5977, 
    287.6157, 287.6355, 287.657, 287.6807, 287.707, 287.7361, 287.4922, 
    287.1841, 286.9031, 286.6455, 286.4084, 286.1899, 285.9875, 285.7996, 
    285.6248, 285.4614, 285.3088, 285.1658, 285.0315, 284.873, 284.6843, 
    284.4958, 284.3074, 284.1187, 283.9302, 283.7417, 283.553, 283.3645, 
    283.176, 282.9875, 282.7988, 282.6104, 282.5938, 282.5771, 282.5608, 
    282.5442, 282.5276, 282.511, 282.4946, 282.478, 282.4614, 282.4448, 
    282.4285, 282.4119, 282.3677, 282.2957, 282.2239, 282.1519, 282.0801, 
    282.0081, 281.936, 281.8643, 281.7922, 281.7205, 281.6484, 281.5767, 
    281.5046, 281.5005, 281.4966, 281.4924, 281.4883, 281.4844, 281.4802, 
    281.4761, 281.4722, 281.468, 281.4639, 281.46, 281.4558, 281.4419, 
    281.4177, 281.3936, 281.3696, 281.3455, 281.3215, 281.2974, 281.2732, 
    281.2493, 281.2251, 281.2012, 281.177, 281.1528, 281.0691, 280.9854, 
    280.9019, 280.8181, 280.7344, 280.6506, 280.5669, 280.4832, 280.3994, 
    280.3157, 280.2319, 280.1482, 280.095, 280.0725, 280.05, 280.0276, 
    280.0051, 279.9827, 279.9602, 279.9377, 279.9153, 279.8928, 279.8704, 
    279.8479, 279.8254, 279.7236, 279.6218, 279.5203, 279.4185, 279.3167, 
    279.2148, 279.113, 279.0115, 278.9097, 278.8079, 278.7061, 278.6045, 
    278.5703, 278.6038, 278.6372, 278.6707, 278.7041, 278.7378, 278.7712, 
    278.8047, 278.8381, 278.8716, 278.905, 278.9385, 278.9722,
  287.1306, 287.1809, 287.231, 287.2812, 287.3315, 287.3816, 287.4319, 
    287.4822, 287.5322, 287.5825, 287.6326, 287.675, 287.7175, 287.76, 
    287.8025, 287.8447, 287.8872, 287.9297, 287.9722, 288.0144, 288.0569, 
    288.0994, 288.1418, 288.1707, 288.186, 288.2014, 288.2168, 288.2322, 
    288.2473, 288.2627, 288.2781, 288.2935, 288.3088, 288.3242, 288.3396, 
    288.355, 288.3364, 288.3181, 288.2996, 288.2812, 288.2627, 288.2444, 
    288.2258, 288.2075, 288.189, 288.1707, 288.1521, 288.1338, 288.1343, 
    288.1538, 288.1733, 288.1929, 288.2124, 288.2319, 288.2515, 288.271, 
    288.2905, 288.3101, 288.3296, 288.3491, 288.3687, 288.3467, 288.3247, 
    288.3025, 288.2805, 288.2585, 288.2363, 288.2144, 288.1921, 288.1702, 
    288.1482, 288.126, 288.104, 288.0713, 288.0283, 287.9851, 287.9419, 
    287.8989, 287.8557, 287.8125, 287.7695, 287.7263, 287.6831, 287.6401, 
    287.5969, 287.5537, 287.5581, 287.5623, 287.5667, 287.5708, 287.5752, 
    287.5793, 287.5837, 287.5879, 287.5923, 287.5964, 287.6008, 287.605, 
    287.5984, 287.5808, 287.5635, 287.5459, 287.5283, 287.5107, 287.4934, 
    287.4758, 287.4583, 287.4409, 287.4233, 287.4058, 287.3882, 287.4084, 
    287.4285, 287.4485, 287.4688, 287.4888, 287.5088, 287.5291, 287.5491, 
    287.5691, 287.5894, 287.6094, 287.6294, 287.6335, 287.6218, 287.6101, 
    287.5984, 287.5867, 287.575, 287.5632, 287.5515, 287.5396, 287.5278, 
    287.5161, 287.5044, 287.4927, 287.4927, 287.4927, 287.4924, 287.4924, 
    287.4924, 287.4924, 287.4924, 287.4924, 287.4922, 287.4922, 287.4922, 
    287.4922, 287.5007, 287.5183, 287.5371, 287.5569, 287.5776, 287.5999, 
    287.623, 287.6479, 287.6743, 287.7024, 287.7324, 287.7644, 287.5291, 
    287.2051, 286.9241, 286.6777, 286.4602, 286.2668, 286.0935, 285.9375, 
    285.7961, 285.6677, 285.5503, 285.4429, 285.3438, 285.1958, 284.9934, 
    284.7908, 284.5884, 284.386, 284.1836, 283.981, 283.7786, 283.5762, 
    283.3735, 283.1711, 282.9688, 282.7661, 282.7339, 282.7014, 282.6689, 
    282.6365, 282.6042, 282.5718, 282.5393, 282.5068, 282.4746, 282.4421, 
    282.4097, 282.3772, 282.3237, 282.2488, 282.1741, 282.0991, 282.0244, 
    281.9495, 281.8748, 281.7998, 281.7251, 281.6501, 281.5754, 281.5005, 
    281.4258, 281.4292, 281.4326, 281.4363, 281.4397, 281.4431, 281.4468, 
    281.4502, 281.4536, 281.4573, 281.4607, 281.4641, 281.4675, 281.4526, 
    281.4194, 281.3862, 281.3528, 281.3196, 281.2861, 281.2529, 281.2197, 
    281.1863, 281.1531, 281.1199, 281.0864, 281.0532, 280.9766, 280.8999, 
    280.8235, 280.7468, 280.6702, 280.5935, 280.5171, 280.4404, 280.3638, 
    280.2871, 280.2107, 280.134, 280.0918, 280.084, 280.0759, 280.0681, 
    280.0603, 280.0525, 280.0447, 280.0366, 280.0288, 280.021, 280.0132, 
    280.0054, 279.9973, 279.8762, 279.7551, 279.634, 279.5127, 279.3916, 
    279.2705, 279.1494, 279.0281, 278.907, 278.7859, 278.6648, 278.5435, 
    278.5007, 278.5364, 278.5723, 278.6079, 278.6436, 278.6792, 278.7148, 
    278.7505, 278.7861, 278.822, 278.8577, 278.8933, 278.929,
  287.1973, 287.2463, 287.2954, 287.3445, 287.3933, 287.4424, 287.4915, 
    287.5405, 287.5896, 287.6387, 287.6877, 287.7285, 287.7695, 287.8105, 
    287.8513, 287.8923, 287.9331, 287.9741, 288.0149, 288.0559, 288.0969, 
    288.1377, 288.1787, 288.2065, 288.2217, 288.2366, 288.2517, 288.2666, 
    288.2815, 288.2966, 288.3115, 288.3267, 288.3416, 288.3567, 288.3716, 
    288.3865, 288.3643, 288.3418, 288.3196, 288.2971, 288.2747, 288.2524, 
    288.23, 288.2078, 288.1853, 288.1628, 288.1406, 288.1182, 288.1177, 
    288.1392, 288.1606, 288.1821, 288.2036, 288.2251, 288.2466, 288.2681, 
    288.2896, 288.311, 288.3325, 288.354, 288.3755, 288.3564, 288.3374, 
    288.3186, 288.2996, 288.2805, 288.2615, 288.2427, 288.2236, 288.2046, 
    288.1858, 288.1667, 288.1477, 288.114, 288.0659, 288.0178, 287.9695, 
    287.9214, 287.873, 287.825, 287.7766, 287.7285, 287.6804, 287.6321, 
    287.584, 287.5356, 287.5359, 287.5359, 287.5359, 287.5361, 287.5361, 
    287.5364, 287.5364, 287.5364, 287.5366, 287.5366, 287.5366, 287.5369, 
    287.5303, 287.5171, 287.5039, 287.4907, 287.4775, 287.4644, 287.4512, 
    287.438, 287.4248, 287.4116, 287.3984, 287.3853, 287.3721, 287.3938, 
    287.4153, 287.4368, 287.4583, 287.48, 287.5015, 287.5229, 287.5444, 
    287.5662, 287.5876, 287.6091, 287.6306, 287.635, 287.6218, 287.6086, 
    287.5957, 287.5825, 287.5693, 287.5564, 287.5432, 287.53, 287.5168, 
    287.5039, 287.4907, 287.4775, 287.4766, 287.4753, 287.4744, 287.4731, 
    287.4722, 287.4709, 287.47, 287.4688, 287.4678, 287.4666, 287.4653, 
    287.4644, 287.4753, 287.499, 287.5232, 287.5486, 287.5747, 287.6016, 
    287.6294, 287.6584, 287.6885, 287.7195, 287.752, 287.7854, 287.5872, 
    287.2358, 286.9529, 286.7202, 286.5254, 286.3601, 286.2178, 286.0942, 
    285.9856, 285.8899, 285.8044, 285.7278, 285.6589, 285.5188, 285.3022, 
    285.0859, 284.8696, 284.6531, 284.4368, 284.2205, 284.0042, 283.7876, 
    283.5713, 283.355, 283.1384, 282.9221, 282.8738, 282.8254, 282.7773, 
    282.729, 282.6807, 282.6323, 282.5842, 282.5359, 282.4875, 282.4392, 
    282.3909, 282.3428, 282.2798, 282.2019, 282.1243, 282.0464, 281.9688, 
    281.8909, 281.8132, 281.7356, 281.6577, 281.5801, 281.5022, 281.4246, 
    281.3467, 281.3579, 281.3689, 281.3799, 281.3911, 281.4021, 281.4131, 
    281.4241, 281.4353, 281.4463, 281.4573, 281.4683, 281.4795, 281.4636, 
    281.4211, 281.3787, 281.3362, 281.2937, 281.251, 281.2085, 281.166, 
    281.1235, 281.0811, 281.0386, 280.9958, 280.9534, 280.884, 280.8145, 
    280.7451, 280.6755, 280.6062, 280.5366, 280.4673, 280.3977, 280.3284, 
    280.2588, 280.1892, 280.1199, 280.0886, 280.0952, 280.1021, 280.1086, 
    280.1155, 280.1223, 280.1289, 280.1357, 280.1426, 280.1492, 280.156, 
    280.1626, 280.1694, 280.0288, 279.8884, 279.7478, 279.6072, 279.4666, 
    279.3259, 279.1855, 279.0449, 278.9043, 278.7637, 278.6233, 278.4827, 
    278.4314, 278.4692, 278.5071, 278.5449, 278.5828, 278.6206, 278.6587, 
    278.6965, 278.7344, 278.7722, 278.8101, 278.8481, 278.886,
  287.2639, 287.3118, 287.3596, 287.4075, 287.4553, 287.5032, 287.5513, 
    287.5991, 287.647, 287.6948, 287.7427, 287.7822, 287.8215, 287.8608, 
    287.9004, 287.9397, 287.9792, 288.0186, 288.0579, 288.0974, 288.1367, 
    288.176, 288.2156, 288.2427, 288.2573, 288.2717, 288.2864, 288.301, 
    288.3157, 288.3303, 288.345, 288.3596, 288.3743, 288.3889, 288.4036, 
    288.4182, 288.3918, 288.3657, 288.3394, 288.313, 288.2866, 288.2605, 
    288.2341, 288.2078, 288.1816, 288.1553, 288.1289, 288.1025, 288.1013, 
    288.1245, 288.1479, 288.1714, 288.1948, 288.2183, 288.2417, 288.2651, 
    288.2886, 288.3118, 288.3352, 288.3586, 288.3821, 288.3662, 288.3503, 
    288.3345, 288.3186, 288.3027, 288.2869, 288.271, 288.2551, 288.239, 
    288.2231, 288.2073, 288.1914, 288.157, 288.1035, 288.0503, 287.9971, 
    287.9438, 287.8906, 287.8372, 287.7839, 287.7307, 287.6775, 287.6243, 
    287.5708, 287.5176, 287.5137, 287.5095, 287.5054, 287.5012, 287.4973, 
    287.4932, 287.489, 287.4849, 287.481, 287.4768, 287.4727, 287.4685, 
    287.4622, 287.4534, 287.4446, 287.4355, 287.4268, 287.418, 287.4092, 
    287.4001, 287.3914, 287.3826, 287.3738, 287.365, 287.356, 287.3792, 
    287.4021, 287.425, 287.448, 287.4709, 287.4939, 287.5171, 287.54, 
    287.563, 287.5859, 287.6089, 287.6318, 287.6362, 287.6218, 287.6072, 
    287.5928, 287.5784, 287.564, 287.5493, 287.5349, 287.5205, 287.5061, 
    287.4915, 287.4771, 287.4626, 287.4604, 287.4583, 287.4561, 287.4539, 
    287.4517, 287.4495, 287.4475, 287.4453, 287.4431, 287.4409, 287.4387, 
    287.4365, 287.4502, 287.48, 287.51, 287.5408, 287.5718, 287.6033, 
    287.635, 287.6675, 287.7002, 287.7336, 287.7673, 287.8018, 287.8364, 
    287.8015, 287.7615, 287.7151, 287.6611, 287.5974, 287.521, 287.4275, 
    287.3105, 286.1296, 286.072, 286.0215, 285.9771, 285.8416, 285.6113, 
    285.3811, 285.1506, 284.9204, 284.6902, 284.4597, 284.2295, 283.9993, 
    283.7688, 283.5386, 283.3083, 283.0781, 283.0139, 282.9497, 282.8855, 
    282.8213, 282.7573, 282.6931, 282.6289, 282.5647, 282.5005, 282.4365, 
    282.3723, 282.3081, 282.2356, 282.155, 282.0745, 281.9937, 281.9131, 
    281.8325, 281.7517, 281.6711, 281.5906, 281.5098, 281.4292, 281.3486, 
    281.2678, 281.2864, 281.3052, 281.3237, 281.3423, 281.3608, 281.3796, 
    281.3982, 281.4167, 281.4353, 281.4541, 281.4727, 281.4912, 281.4746, 
    281.4229, 281.3711, 281.3193, 281.2676, 281.2158, 281.1641, 281.1123, 
    281.0605, 281.0088, 280.957, 280.9055, 280.8538, 280.7913, 280.729, 
    280.6667, 280.6042, 280.542, 280.4797, 280.4175, 280.355, 280.2927, 
    280.2305, 280.168, 280.1057, 280.0852, 280.1067, 280.1279, 280.1494, 
    280.1707, 280.1919, 280.2134, 280.2346, 280.2561, 280.2773, 280.2988, 
    280.3201, 280.3416, 280.1814, 280.0215, 279.8616, 279.7017, 279.5415, 
    279.3816, 279.2217, 279.0618, 278.9016, 278.7417, 278.5818, 278.4219, 
    278.3618, 278.4019, 278.4419, 278.4822, 278.5222, 278.5623, 278.6023, 
    278.6423, 278.6826, 278.7227, 278.7627, 278.8027, 278.8428,
  287.3103, 287.3582, 287.406, 287.4539, 287.5017, 287.5496, 287.5974, 
    287.6453, 287.6931, 287.741, 287.7888, 287.8271, 287.8655, 287.9038, 
    287.9421, 287.9805, 288.0188, 288.0571, 288.0952, 288.1335, 288.1719, 
    288.2102, 288.2485, 288.2747, 288.2886, 288.3027, 288.3167, 288.3306, 
    288.3445, 288.3586, 288.3726, 288.3865, 288.4004, 288.4146, 288.4285, 
    288.4424, 288.4141, 288.3855, 288.3572, 288.3286, 288.3003, 288.2717, 
    288.2434, 288.2148, 288.1865, 288.158, 288.1296, 288.1011, 288.0986, 
    288.1223, 288.1458, 288.1692, 288.1929, 288.2163, 288.2397, 288.2634, 
    288.2869, 288.3103, 288.334, 288.3574, 288.3809, 288.3674, 288.354, 
    288.3406, 288.3269, 288.3135, 288.3, 288.2864, 288.2729, 288.2595, 
    288.2458, 288.2324, 288.219, 288.1838, 288.1274, 288.0708, 288.0142, 
    287.9578, 287.9011, 287.8445, 287.7881, 287.7314, 287.6748, 287.6184, 
    287.5618, 287.5051, 287.4978, 287.4905, 287.4832, 287.4758, 287.4685, 
    287.4609, 287.4536, 287.4463, 287.439, 287.4316, 287.4241, 287.4167, 
    287.4104, 287.4048, 287.3992, 287.3936, 287.3879, 287.3823, 287.3767, 
    287.3711, 287.3655, 287.3599, 287.3542, 287.3486, 287.3433, 287.366, 
    287.3884, 287.4111, 287.4338, 287.4565, 287.4792, 287.502, 287.5247, 
    287.5474, 287.5701, 287.5928, 287.6155, 287.6199, 287.6062, 287.5925, 
    287.5789, 287.5652, 287.5515, 287.5378, 287.5242, 287.5105, 287.4968, 
    287.4832, 287.4692, 287.4556, 287.4534, 287.4509, 287.4487, 287.4465, 
    287.4441, 287.4419, 287.4395, 287.4373, 287.4348, 287.4326, 287.4302, 
    287.428, 287.4431, 287.4756, 287.5081, 287.5405, 287.5732, 287.6057, 
    287.6382, 287.6707, 287.7031, 287.7358, 287.7683, 287.8008, 287.8333, 
    287.8044, 287.7712, 287.7329, 287.688, 287.6345, 287.5701, 287.4905, 
    287.3901, 286.2659, 286.2244, 286.1887, 286.1577, 286.0234, 285.7825, 
    285.5417, 285.3008, 285.0598, 284.8191, 284.5781, 284.3372, 284.0964, 
    283.8555, 283.6145, 283.3738, 283.1328, 283.0605, 282.9885, 282.9163, 
    282.844, 282.772, 282.6997, 282.6274, 282.5552, 282.4832, 282.4109, 
    282.3386, 282.2666, 282.1897, 282.1079, 282.0264, 281.9446, 281.863, 
    281.7812, 281.6997, 281.6182, 281.5364, 281.4548, 281.373, 281.2915, 
    281.2097, 281.2317, 281.2534, 281.2754, 281.2971, 281.3191, 281.3408, 
    281.3625, 281.3845, 281.4062, 281.4282, 281.45, 281.4719, 281.4541, 
    281.3967, 281.3396, 281.2822, 281.2251, 281.1677, 281.1106, 281.0532, 
    280.9961, 280.9387, 280.8816, 280.8242, 280.7671, 280.7104, 280.6541, 
    280.5974, 280.541, 280.4844, 280.428, 280.3713, 280.3149, 280.2585, 
    280.2019, 280.1455, 280.0889, 280.075, 280.1035, 280.1321, 280.1606, 
    280.1892, 280.2178, 280.2463, 280.2749, 280.3035, 280.3323, 280.3608, 
    280.3894, 280.418, 280.2478, 280.0779, 279.908, 279.7378, 279.5679, 
    279.3977, 279.2278, 279.0579, 278.8877, 278.7178, 278.5476, 278.3777, 
    278.3135, 278.3552, 278.397, 278.4387, 278.4805, 278.5222, 278.564, 
    278.6057, 278.6475, 278.6892, 278.731, 278.7727, 278.8145,
  287.2986, 287.3496, 287.4006, 287.4519, 287.5029, 287.554, 287.605, 
    287.6562, 287.7073, 287.7583, 287.8093, 287.8479, 287.8862, 287.9246, 
    287.9631, 288.0015, 288.04, 288.0784, 288.1167, 288.1553, 288.1936, 
    288.2319, 288.2705, 288.2959, 288.3083, 288.3208, 288.3333, 288.3455, 
    288.3579, 288.3704, 288.3828, 288.3953, 288.4077, 288.4202, 288.4324, 
    288.4448, 288.4194, 288.394, 288.3687, 288.3433, 288.3179, 288.2925, 
    288.2671, 288.2417, 288.2163, 288.1909, 288.1655, 288.1401, 288.1367, 
    288.155, 288.1736, 288.1919, 288.2102, 288.2288, 288.2471, 288.2654, 
    288.2837, 288.3022, 288.3206, 288.3389, 288.3574, 288.3442, 288.3311, 
    288.3179, 288.3047, 288.2915, 288.2786, 288.2654, 288.2522, 288.239, 
    288.2258, 288.2126, 288.1995, 288.1658, 288.1108, 288.0562, 288.0015, 
    287.9468, 287.8921, 287.8374, 287.7827, 287.728, 287.6733, 287.6187, 
    287.564, 287.509, 287.501, 287.4929, 287.4849, 287.4768, 287.4688, 
    287.4607, 287.4526, 287.4446, 287.4363, 287.4282, 287.4202, 287.4121, 
    287.4053, 287.3999, 287.3943, 287.3889, 287.3833, 287.3779, 287.3726, 
    287.3669, 287.3616, 287.356, 287.3506, 287.345, 287.3396, 287.3569, 
    287.3743, 287.3916, 287.4089, 287.4265, 287.4438, 287.4612, 287.4785, 
    287.4958, 287.5134, 287.5308, 287.5481, 287.5535, 287.5466, 287.5398, 
    287.533, 287.5261, 287.5193, 287.5127, 287.5059, 287.499, 287.4922, 
    287.4854, 287.4785, 287.4717, 287.4719, 287.4722, 287.4724, 287.4727, 
    287.4729, 287.4734, 287.4736, 287.4739, 287.4741, 287.4744, 287.4746, 
    287.4749, 287.4873, 287.512, 287.5366, 287.5613, 287.5862, 287.6108, 
    287.6355, 287.6602, 287.6851, 287.7097, 287.7344, 287.759, 287.7837, 
    287.752, 287.7153, 287.6731, 287.6235, 287.5647, 287.4934, 287.4058, 
    287.2952, 286.0549, 286.0093, 285.97, 285.9358, 285.7996, 285.5576, 
    285.3157, 285.0737, 284.832, 284.5901, 284.3481, 284.1062, 283.8645, 
    283.6226, 283.3806, 283.1387, 282.897, 282.8391, 282.7815, 282.7239, 
    282.6663, 282.6086, 282.5508, 282.4932, 282.4355, 282.3779, 282.3201, 
    282.2625, 282.2048, 282.1375, 282.0603, 281.9832, 281.906, 281.8289, 
    281.7517, 281.6746, 281.5974, 281.5203, 281.4431, 281.366, 281.2888, 
    281.2117, 281.2244, 281.2368, 281.2495, 281.2622, 281.2747, 281.2874, 
    281.2998, 281.3125, 281.325, 281.3376, 281.3501, 281.3628, 281.343, 
    281.291, 281.2388, 281.1868, 281.1348, 281.0828, 281.0305, 280.9785, 
    280.9265, 280.8743, 280.8223, 280.7703, 280.718, 280.6636, 280.6091, 
    280.5547, 280.5002, 280.4456, 280.3911, 280.3367, 280.2822, 280.2278, 
    280.1733, 280.1187, 280.0642, 280.0444, 280.0588, 280.0735, 280.0881, 
    280.1028, 280.1172, 280.1318, 280.1465, 280.1611, 280.1758, 280.1902, 
    280.2048, 280.2195, 280.0664, 279.9133, 279.76, 279.6069, 279.4539, 
    279.3008, 279.1477, 278.9946, 278.8413, 278.6882, 278.5352, 278.3821, 
    278.3264, 278.3682, 278.4102, 278.4519, 278.4939, 278.5356, 278.5776, 
    278.6194, 278.6614, 278.7031, 278.7449, 278.7869, 278.8286,
  287.2869, 287.3411, 287.3955, 287.4497, 287.5042, 287.5583, 287.6128, 
    287.667, 287.7214, 287.7756, 287.8301, 287.8684, 287.907, 287.9456, 
    287.9841, 288.0227, 288.0613, 288.0996, 288.1382, 288.1768, 288.2153, 
    288.2539, 288.2922, 288.3171, 288.3279, 288.3389, 288.3496, 288.3606, 
    288.3713, 288.3823, 288.3931, 288.4041, 288.4148, 288.4258, 288.4365, 
    288.4475, 288.425, 288.4026, 288.3804, 288.3579, 288.3357, 288.3132, 
    288.291, 288.2686, 288.2463, 288.2239, 288.2017, 288.1792, 288.1748, 
    288.188, 288.2012, 288.2146, 288.2278, 288.241, 288.2542, 288.2676, 
    288.2808, 288.2939, 288.3071, 288.3206, 288.3337, 288.321, 288.3081, 
    288.2954, 288.2825, 288.2698, 288.2571, 288.2441, 288.2314, 288.2185, 
    288.2058, 288.1931, 288.1802, 288.1475, 288.0945, 288.0417, 287.9888, 
    287.936, 287.8831, 287.8303, 287.7773, 287.7244, 287.6716, 287.6187, 
    287.5659, 287.5129, 287.5042, 287.4954, 287.4866, 287.4778, 287.469, 
    287.4602, 287.4514, 287.4426, 287.4338, 287.425, 287.4163, 287.4075, 
    287.4004, 287.395, 287.3896, 287.3843, 287.3789, 287.3735, 287.3682, 
    287.3628, 287.3574, 287.3521, 287.3467, 287.3413, 287.3359, 287.3479, 
    287.3601, 287.3721, 287.3843, 287.3962, 287.4082, 287.4204, 287.4324, 
    287.4446, 287.4565, 287.4688, 287.4807, 287.4868, 287.4868, 287.4871, 
    287.4871, 287.4871, 287.4873, 287.4873, 287.4875, 287.4875, 287.4875, 
    287.4878, 287.4878, 287.4878, 287.4907, 287.4934, 287.4963, 287.499, 
    287.502, 287.5046, 287.5076, 287.5103, 287.5132, 287.5159, 287.5188, 
    287.5215, 287.5315, 287.5483, 287.5652, 287.582, 287.5991, 287.616, 
    287.6328, 287.6499, 287.6667, 287.6836, 287.7004, 287.7175, 287.7344, 
    287.6995, 287.6597, 287.6133, 287.5591, 287.4946, 287.4167, 287.321, 
    287.2, 285.844, 285.7939, 285.7512, 285.7139, 285.5757, 285.3328, 
    285.0898, 284.8469, 284.604, 284.3611, 284.1182, 283.8755, 283.6326, 
    283.3896, 283.1467, 282.9038, 282.6609, 282.6179, 282.5747, 282.5315, 
    282.4883, 282.4451, 282.4021, 282.3589, 282.3157, 282.2725, 282.2295, 
    282.1863, 282.1431, 282.0852, 282.0125, 281.9399, 281.8674, 281.7947, 
    281.7222, 281.6494, 281.5769, 281.5042, 281.4316, 281.3589, 281.2864, 
    281.2136, 281.217, 281.2205, 281.2236, 281.2271, 281.2305, 281.2336, 
    281.2371, 281.2405, 281.2437, 281.2471, 281.2505, 281.2537, 281.2319, 
    281.1851, 281.1382, 281.0913, 281.0444, 280.9976, 280.9507, 280.9038, 
    280.8567, 280.8098, 280.7629, 280.7161, 280.6692, 280.6167, 280.5642, 
    280.5117, 280.4592, 280.407, 280.3545, 280.302, 280.2495, 280.197, 
    280.1445, 280.092, 280.0396, 280.0137, 280.0144, 280.0149, 280.0156, 
    280.0161, 280.0168, 280.0173, 280.0181, 280.0186, 280.0193, 280.0198, 
    280.0205, 280.021, 279.8848, 279.7485, 279.6123, 279.4761, 279.3398, 
    279.2036, 279.0674, 278.9312, 278.7952, 278.6589, 278.5227, 278.3865, 
    278.3394, 278.3811, 278.4231, 278.4651, 278.5071, 278.5491, 278.5911, 
    278.6331, 278.675, 278.717, 278.759, 278.801, 278.8428,
  287.2751, 287.3328, 287.3904, 287.4478, 287.5054, 287.563, 287.6204, 
    287.678, 287.7354, 287.793, 287.8506, 287.8892, 287.9277, 287.9666, 
    288.0051, 288.0437, 288.0823, 288.1211, 288.1597, 288.1982, 288.2371, 
    288.2756, 288.3142, 288.3381, 288.3477, 288.3569, 288.3662, 288.3755, 
    288.3848, 288.394, 288.4033, 288.4126, 288.4219, 288.4314, 288.4407, 
    288.45, 288.4307, 288.4114, 288.3921, 288.3728, 288.3535, 288.3342, 
    288.3147, 288.2954, 288.2761, 288.2568, 288.2375, 288.2183, 288.2126, 
    288.2209, 288.229, 288.2371, 288.2451, 288.2534, 288.2615, 288.2695, 
    288.2776, 288.2856, 288.2939, 288.302, 288.3101, 288.2976, 288.2852, 
    288.2727, 288.2603, 288.248, 288.2356, 288.2231, 288.2107, 288.1982, 
    288.1858, 288.1733, 288.1609, 288.1292, 288.0781, 288.0271, 287.9761, 
    287.925, 287.874, 287.823, 287.772, 287.7209, 287.6699, 287.6189, 
    287.5679, 287.5168, 287.5073, 287.4978, 287.4883, 287.479, 287.4695, 
    287.46, 287.4504, 287.4409, 287.4314, 287.4219, 287.4124, 287.4028, 
    287.3955, 287.3901, 287.385, 287.3796, 287.3745, 287.3691, 287.364, 
    287.3586, 287.3533, 287.3481, 287.3428, 287.3376, 287.3323, 287.3391, 
    287.3457, 287.3525, 287.3594, 287.366, 287.3728, 287.3796, 287.3862, 
    287.3931, 287.3999, 287.4065, 287.4133, 287.4202, 287.4272, 287.4341, 
    287.4412, 287.4482, 287.4551, 287.4622, 287.469, 287.4761, 287.4832, 
    287.49, 287.4971, 287.5039, 287.5093, 287.5146, 287.52, 287.5254, 
    287.5308, 287.5361, 287.5415, 287.5469, 287.5522, 287.5576, 287.563, 
    287.5684, 287.5757, 287.5847, 287.5938, 287.603, 287.6121, 287.6211, 
    287.6301, 287.6394, 287.6484, 287.6575, 287.6667, 287.6758, 287.6848, 
    287.647, 287.6038, 287.5535, 287.4946, 287.4248, 287.3403, 287.2363, 
    287.105, 285.6333, 285.5789, 285.5322, 285.4919, 285.3516, 285.1077, 
    284.864, 284.6201, 284.3762, 284.1323, 283.8884, 283.6445, 283.4006, 
    283.1567, 282.9128, 282.6689, 282.425, 282.3965, 282.3677, 282.3391, 
    282.3105, 282.2817, 282.2532, 282.2246, 282.1958, 282.1672, 282.1387, 
    282.1101, 282.0813, 282.033, 281.9648, 281.8967, 281.8286, 281.7605, 
    281.6924, 281.6243, 281.5562, 281.488, 281.4199, 281.3518, 281.2837, 
    281.2156, 281.2097, 281.2039, 281.198, 281.1919, 281.186, 281.1802, 
    281.1743, 281.1685, 281.1624, 281.1565, 281.1506, 281.1448, 281.1208, 
    281.0791, 281.0374, 280.9958, 280.9541, 280.9124, 280.8706, 280.8289, 
    280.7871, 280.7454, 280.7036, 280.6621, 280.6204, 280.5698, 280.5195, 
    280.469, 280.4185, 280.3682, 280.3176, 280.2671, 280.2168, 280.1663, 
    280.116, 280.0654, 280.0149, 279.9832, 279.9697, 279.9563, 279.9429, 
    279.9297, 279.9163, 279.9028, 279.8894, 279.8762, 279.8628, 279.8494, 
    279.8359, 279.8228, 279.7034, 279.584, 279.4646, 279.3455, 279.2261, 
    279.1067, 278.9873, 278.8679, 278.7488, 278.6294, 278.51, 278.3906, 
    278.3521, 278.3943, 278.4363, 278.4783, 278.5205, 278.5625, 278.6045, 
    278.6467, 278.6887, 278.7307, 278.7729, 278.8149, 278.8569,
  287.2634, 287.3242, 287.385, 287.4458, 287.5066, 287.5674, 287.6282, 
    287.6887, 287.7495, 287.8103, 287.8711, 287.9099, 287.9485, 287.9873, 
    288.0261, 288.0649, 288.1035, 288.1423, 288.1812, 288.22, 288.2585, 
    288.2974, 288.3362, 288.3594, 288.3672, 288.375, 288.3826, 288.3904, 
    288.3982, 288.406, 288.4136, 288.4214, 288.4292, 288.437, 288.4446, 
    288.4524, 288.436, 288.4199, 288.4036, 288.3875, 288.3711, 288.355, 
    288.3386, 288.3223, 288.3062, 288.2898, 288.2737, 288.2573, 288.2507, 
    288.2537, 288.2566, 288.2598, 288.2627, 288.2656, 288.2686, 288.2715, 
    288.2747, 288.2776, 288.2805, 288.2834, 288.2864, 288.2744, 288.2622, 
    288.2502, 288.2383, 288.2261, 288.2141, 288.2019, 288.1899, 288.1777, 
    288.1658, 288.1536, 288.1416, 288.1108, 288.0618, 288.0125, 287.9634, 
    287.9143, 287.865, 287.8159, 287.7666, 287.7175, 287.6682, 287.6191, 
    287.5701, 287.5208, 287.5105, 287.5005, 287.4902, 287.48, 287.4697, 
    287.4595, 287.4492, 287.439, 287.429, 287.4187, 287.4084, 287.3982, 
    287.3906, 287.3853, 287.3801, 287.375, 287.3699, 287.3647, 287.3596, 
    287.3545, 287.3494, 287.3442, 287.3391, 287.3337, 287.3286, 287.3301, 
    287.3315, 287.333, 287.3345, 287.3359, 287.3374, 287.3389, 287.3403, 
    287.3416, 287.343, 287.3445, 287.3459, 287.3535, 287.3674, 287.3813, 
    287.3953, 287.4092, 287.4231, 287.4368, 287.4507, 287.4646, 287.4785, 
    287.4924, 287.5063, 287.52, 287.5281, 287.5359, 287.5439, 287.5518, 
    287.5598, 287.5676, 287.5754, 287.5835, 287.5913, 287.5994, 287.6072, 
    287.6152, 287.6199, 287.6211, 287.6223, 287.6238, 287.625, 287.6262, 
    287.6277, 287.6289, 287.6301, 287.6316, 287.6328, 287.634, 287.6355, 
    287.5947, 287.5479, 287.4937, 287.4302, 287.3547, 287.2637, 287.1514, 
    287.0098, 285.4224, 285.3638, 285.3135, 285.2698, 285.1277, 284.8828, 
    284.6379, 284.3931, 284.1482, 283.9033, 283.6584, 283.4136, 283.1687, 
    282.9238, 282.679, 282.4341, 282.1892, 282.175, 282.1609, 282.1467, 
    282.1326, 282.1184, 282.1045, 282.0903, 282.0762, 282.062, 282.0479, 
    282.0337, 282.0195, 281.9807, 281.9172, 281.8535, 281.79, 281.7263, 
    281.6628, 281.5991, 281.5356, 281.4719, 281.4084, 281.3447, 281.2812, 
    281.2175, 281.2024, 281.1873, 281.1721, 281.157, 281.1418, 281.1267, 
    281.1116, 281.0964, 281.0811, 281.0659, 281.0508, 281.0356, 281.0098, 
    280.9734, 280.9368, 280.9001, 280.8638, 280.8271, 280.7905, 280.7542, 
    280.7175, 280.6809, 280.6445, 280.6079, 280.5713, 280.5229, 280.4746, 
    280.426, 280.3777, 280.3293, 280.2808, 280.2324, 280.1841, 280.1357, 
    280.0872, 280.0388, 279.9905, 279.9524, 279.925, 279.8977, 279.8704, 
    279.843, 279.8157, 279.7883, 279.761, 279.7336, 279.7063, 279.679, 
    279.6516, 279.6243, 279.5217, 279.4194, 279.3169, 279.2146, 279.1121, 
    279.0098, 278.9072, 278.8047, 278.7024, 278.5999, 278.4976, 278.395, 
    278.365, 278.4072, 278.4492, 278.4915, 278.5337, 278.5759, 278.6182, 
    278.6602, 278.7024, 278.7446, 278.7869, 278.8291, 278.8713,
  287.252, 287.3159, 287.3799, 287.4438, 287.5078, 287.5718, 287.6357, 
    287.6997, 287.7637, 287.8276, 287.8916, 287.9304, 287.9695, 288.0083, 
    288.0471, 288.0859, 288.1248, 288.1638, 288.2026, 288.2415, 288.2803, 
    288.3191, 288.3582, 288.3806, 288.3867, 288.3931, 288.3992, 288.4053, 
    288.4116, 288.4177, 288.4238, 288.4302, 288.4363, 288.4426, 288.4487, 
    288.4548, 288.4417, 288.4285, 288.4153, 288.4021, 288.3889, 288.3757, 
    288.3625, 288.3494, 288.3359, 288.3228, 288.3096, 288.2964, 288.2888, 
    288.2866, 288.2844, 288.2822, 288.28, 288.2781, 288.2759, 288.2737, 
    288.2715, 288.2693, 288.2671, 288.2651, 288.2629, 288.2512, 288.2395, 
    288.2278, 288.2161, 288.2043, 288.1926, 288.1809, 288.1692, 288.1572, 
    288.1455, 288.1338, 288.1221, 288.0925, 288.0454, 287.998, 287.9507, 
    287.9033, 287.856, 287.8086, 287.7612, 287.7141, 287.6667, 287.6194, 
    287.572, 287.5247, 287.5137, 287.5029, 287.4919, 287.481, 287.47, 
    287.4592, 287.4482, 287.4373, 287.4263, 287.4155, 287.4045, 287.3936, 
    287.3855, 287.3806, 287.3755, 287.3704, 287.3655, 287.3604, 287.3552, 
    287.3503, 287.3452, 287.3403, 287.3352, 287.3301, 287.3252, 287.3213, 
    287.3174, 287.3135, 287.3096, 287.3057, 287.3018, 287.2979, 287.2942, 
    287.2903, 287.2864, 287.2825, 287.2786, 287.2871, 287.3079, 287.3286, 
    287.3494, 287.3701, 287.3909, 287.4116, 287.4324, 287.4531, 287.4739, 
    287.4946, 287.5154, 287.5361, 287.5466, 287.5571, 287.5676, 287.5781, 
    287.5886, 287.5991, 287.6096, 287.6201, 287.6306, 287.6409, 287.6514, 
    287.6619, 287.6638, 287.6575, 287.6509, 287.6445, 287.6379, 287.6313, 
    287.625, 287.6184, 287.6121, 287.6055, 287.5989, 287.5925, 287.5859, 
    287.5422, 287.4919, 287.4338, 287.3657, 287.2849, 287.187, 287.0667, 
    286.9148, 285.2114, 285.1487, 285.0947, 285.0479, 284.9038, 284.658, 
    284.4121, 284.1663, 283.9202, 283.6743, 283.4285, 283.1826, 282.9368, 
    282.6909, 282.4451, 282.199, 281.9531, 281.9536, 281.9541, 281.9543, 
    281.9548, 281.9551, 281.9556, 281.9561, 281.9563, 281.9568, 281.957, 
    281.9575, 281.958, 281.9285, 281.8694, 281.8103, 281.7512, 281.6921, 
    281.6331, 281.574, 281.5149, 281.4558, 281.3967, 281.3376, 281.2786, 
    281.2195, 281.1951, 281.1707, 281.1462, 281.1218, 281.0974, 281.073, 
    281.0486, 281.0242, 281, 280.9756, 280.9512, 280.9268, 280.8987, 
    280.8674, 280.8359, 280.8047, 280.7734, 280.7419, 280.7107, 280.6792, 
    280.6479, 280.6165, 280.5852, 280.5537, 280.5225, 280.4761, 280.4297, 
    280.3833, 280.3369, 280.2905, 280.2441, 280.1978, 280.1514, 280.105, 
    280.0586, 280.0122, 279.9658, 279.9219, 279.8806, 279.8391, 279.7979, 
    279.7566, 279.7151, 279.6738, 279.6326, 279.5913, 279.5498, 279.5085, 
    279.4673, 279.4258, 279.3403, 279.2549, 279.1692, 279.0837, 278.998, 
    278.9126, 278.8271, 278.7415, 278.656, 278.5706, 278.4849, 278.3994, 
    278.3777, 278.4202, 278.4624, 278.5046, 278.5469, 278.5894, 278.6316, 
    278.6738, 278.7163, 278.7585, 278.8008, 278.843, 278.8855,
  287.2402, 287.3074, 287.3745, 287.4419, 287.509, 287.5762, 287.6433, 
    287.7107, 287.7778, 287.845, 287.9121, 287.9512, 287.9902, 288.0291, 
    288.0681, 288.1072, 288.146, 288.1851, 288.2241, 288.2629, 288.302, 
    288.3411, 288.3799, 288.4019, 288.4065, 288.4111, 288.4158, 288.4204, 
    288.425, 288.4297, 288.4343, 288.439, 288.4436, 288.448, 288.4526, 
    288.4573, 288.4473, 288.437, 288.427, 288.4167, 288.4065, 288.3965, 
    288.3862, 288.3762, 288.366, 288.3557, 288.3457, 288.3354, 288.3267, 
    288.3196, 288.3123, 288.3049, 288.2976, 288.2903, 288.283, 288.2756, 
    288.2683, 288.2612, 288.2539, 288.2466, 288.2393, 288.2278, 288.2166, 
    288.2051, 288.1938, 288.1824, 288.1711, 288.1597, 288.1482, 288.137, 
    288.1255, 288.1143, 288.1028, 288.0745, 288.0288, 287.9834, 287.938, 
    287.8926, 287.8469, 287.8015, 287.7561, 287.7104, 287.665, 287.6196, 
    287.574, 287.5286, 287.5168, 287.5054, 287.4937, 287.4819, 287.4705, 
    287.4587, 287.447, 287.4355, 287.4238, 287.4121, 287.4006, 287.3889, 
    287.3806, 287.3757, 287.3708, 287.3657, 287.3608, 287.356, 287.3511, 
    287.3462, 287.3413, 287.3362, 287.3313, 287.3264, 287.3215, 287.3123, 
    287.3032, 287.2939, 287.2847, 287.2756, 287.2664, 287.2571, 287.248, 
    287.2388, 287.2295, 287.2205, 287.2112, 287.2205, 287.248, 287.2759, 
    287.3035, 287.3311, 287.3586, 287.3865, 287.4141, 287.4417, 287.4695, 
    287.4971, 287.5247, 287.5525, 287.5654, 287.5784, 287.5916, 287.6045, 
    287.6174, 287.6306, 287.6436, 287.6565, 287.6697, 287.6826, 287.6958, 
    287.7087, 287.708, 287.6938, 287.6794, 287.6653, 287.6509, 287.6365, 
    287.6223, 287.6079, 287.5938, 287.5793, 287.5652, 287.5508, 287.5364, 
    287.4897, 287.4363, 287.374, 287.3013, 287.2148, 287.1106, 286.9819, 
    286.8196, 285.0005, 284.9336, 284.876, 284.8259, 284.6799, 284.4331, 
    284.186, 283.9392, 283.6924, 283.4456, 283.1985, 282.9517, 282.7048, 
    282.458, 282.2109, 281.9641, 281.7173, 281.7322, 281.7471, 281.762, 
    281.7769, 281.7917, 281.8066, 281.8215, 281.8364, 281.8516, 281.8665, 
    281.8813, 281.8962, 281.8765, 281.8218, 281.7671, 281.7126, 281.658, 
    281.6035, 281.5488, 281.4944, 281.4397, 281.3853, 281.3306, 281.2761, 
    281.2214, 281.1877, 281.1543, 281.1206, 281.0869, 281.0532, 281.0195, 
    280.9858, 280.9521, 280.9187, 280.885, 280.8513, 280.8176, 280.7876, 
    280.7615, 280.7354, 280.7092, 280.6831, 280.6567, 280.6306, 280.6045, 
    280.5784, 280.552, 280.5259, 280.4998, 280.4736, 280.4292, 280.3848, 
    280.3403, 280.2961, 280.2517, 280.2073, 280.1631, 280.1187, 280.0742, 
    280.0298, 279.9856, 279.9412, 279.8914, 279.8359, 279.7805, 279.7253, 
    279.6699, 279.6147, 279.5593, 279.5042, 279.4487, 279.3933, 279.3381, 
    279.2827, 279.2275, 279.1587, 279.0901, 279.0215, 278.9529, 278.8843, 
    278.8157, 278.7468, 278.6782, 278.6096, 278.541, 278.4724, 278.4038, 
    278.3906, 278.4331, 278.4753, 278.5178, 278.5603, 278.6028, 278.645, 
    278.6875, 278.73, 278.7722, 278.8147, 278.8572, 278.8997,
  287.2119, 287.2817, 287.3516, 287.4214, 287.4912, 287.561, 287.6309, 
    287.7007, 287.7705, 287.8403, 287.9099, 287.9495, 287.989, 288.0286, 
    288.0681, 288.1077, 288.1472, 288.1865, 288.2261, 288.2656, 288.3052, 
    288.3447, 288.3843, 288.4058, 288.4094, 288.4133, 288.417, 288.4207, 
    288.4243, 288.428, 288.4319, 288.4355, 288.4392, 288.4429, 288.4465, 
    288.4504, 288.4429, 288.4353, 288.4277, 288.4202, 288.4126, 288.405, 
    288.3975, 288.3901, 288.3826, 288.375, 288.3674, 288.3599, 288.3506, 
    288.3398, 288.3289, 288.3179, 288.3069, 288.2961, 288.2852, 288.2742, 
    288.2634, 288.2524, 288.2415, 288.2305, 288.2197, 288.2092, 288.199, 
    288.1887, 288.1785, 288.1682, 288.158, 288.1477, 288.1375, 288.127, 
    288.1167, 288.1064, 288.0962, 288.0686, 288.0239, 287.9792, 287.9348, 
    287.8901, 287.8455, 287.8008, 287.7561, 287.7114, 287.6667, 287.6221, 
    287.5774, 287.5327, 287.52, 287.5076, 287.4949, 287.4824, 287.4697, 
    287.4573, 287.4446, 287.4321, 287.4194, 287.407, 287.3943, 287.3818, 
    287.3735, 287.3694, 287.3655, 287.3613, 287.3574, 287.3533, 287.3494, 
    287.3452, 287.3413, 287.3372, 287.3333, 287.3291, 287.3252, 287.3113, 
    287.2976, 287.2839, 287.27, 287.2563, 287.2427, 287.2288, 287.2151, 
    287.2014, 287.1877, 287.1738, 287.1602, 287.1699, 287.2034, 287.2368, 
    287.2703, 287.3035, 287.3369, 287.3704, 287.4038, 287.4373, 287.4707, 
    287.5042, 287.5374, 287.5708, 287.5857, 287.6006, 287.6157, 287.6306, 
    287.6455, 287.6604, 287.6753, 287.6902, 287.7051, 287.72, 287.7351, 
    287.75, 287.748, 287.729, 287.7102, 287.6912, 287.6724, 287.6533, 
    287.6345, 287.6155, 287.5967, 287.5776, 287.5588, 287.5398, 287.521, 
    287.4729, 287.4177, 287.3538, 287.2791, 287.1899, 287.0825, 286.9502, 
    286.7832, 284.9109, 284.842, 284.7827, 284.7312, 284.5808, 284.3262, 
    284.0715, 283.8171, 283.5625, 283.3081, 283.0535, 282.7991, 282.5444, 
    282.2898, 282.0354, 281.7808, 281.5264, 281.5522, 281.5779, 281.6038, 
    281.6296, 281.6555, 281.6814, 281.7073, 281.7329, 281.7588, 281.7847, 
    281.8105, 281.8364, 281.824, 281.7732, 281.7224, 281.6719, 281.6211, 
    281.5703, 281.5195, 281.469, 281.4182, 281.3674, 281.3167, 281.2661, 
    281.2153, 281.1746, 281.1338, 281.0933, 281.0525, 281.0117, 280.9712, 
    280.9304, 280.8896, 280.8491, 280.8083, 280.7676, 280.7271, 280.6953, 
    280.6729, 280.6504, 280.6279, 280.6055, 280.583, 280.5603, 280.5378, 
    280.5154, 280.4929, 280.4705, 280.448, 280.4255, 280.3828, 280.3403, 
    280.2976, 280.2551, 280.2124, 280.1699, 280.1272, 280.0847, 280.0422, 
    279.9995, 279.957, 279.9143, 279.8601, 279.7944, 279.7288, 279.6631, 
    279.5974, 279.5317, 279.4661, 279.4004, 279.3345, 279.2688, 279.2031, 
    279.1375, 279.0718, 279.0164, 278.9612, 278.9058, 278.8503, 278.7952, 
    278.7397, 278.6846, 278.6292, 278.5737, 278.5186, 278.4631, 278.408, 
    278.4004, 278.4407, 278.481, 278.5212, 278.5615, 278.6018, 278.6421, 
    278.6824, 278.7227, 278.7629, 278.803, 278.8433, 278.8835,
  287.1279, 287.1982, 287.2686, 287.3389, 287.4094, 287.4797, 287.55, 
    287.6204, 287.6907, 287.761, 287.8313, 287.8728, 287.9143, 287.9558, 
    287.9973, 288.0388, 288.0803, 288.1218, 288.1633, 288.2048, 288.2463, 
    288.2878, 288.3293, 288.3525, 288.3574, 288.3623, 288.3672, 288.3721, 
    288.377, 288.3818, 288.3867, 288.3916, 288.3965, 288.4014, 288.4062, 
    288.4111, 288.4048, 288.3984, 288.3921, 288.3857, 288.3794, 288.373, 
    288.3667, 288.3604, 288.354, 288.3479, 288.3416, 288.3352, 288.3271, 
    288.3176, 288.3083, 288.2988, 288.2893, 288.2798, 288.2703, 288.261, 
    288.2515, 288.2419, 288.2324, 288.2229, 288.2136, 288.2068, 288.2, 
    288.1931, 288.1865, 288.1797, 288.1729, 288.166, 288.1594, 288.1526, 
    288.1458, 288.1389, 288.1323, 288.1052, 288.0579, 288.0105, 287.9631, 
    287.916, 287.8687, 287.8213, 287.7739, 287.7266, 287.6794, 287.6321, 
    287.5847, 287.5374, 287.5232, 287.5088, 287.4946, 287.4802, 287.4661, 
    287.4519, 287.4375, 287.4233, 287.4089, 287.3948, 287.3804, 287.3662, 
    287.3589, 287.3584, 287.3579, 287.3574, 287.3569, 287.3564, 287.356, 
    287.3555, 287.355, 287.3545, 287.3542, 287.3538, 287.3533, 287.3374, 
    287.3215, 287.3059, 287.29, 287.2742, 287.2585, 287.2427, 287.2268, 
    287.2109, 287.1953, 287.1794, 287.1636, 287.1733, 287.2087, 287.2441, 
    287.2793, 287.3147, 287.3501, 287.3853, 287.4207, 287.4561, 287.4912, 
    287.5266, 287.562, 287.5972, 287.6118, 287.6265, 287.6411, 287.6555, 
    287.6702, 287.6848, 287.6995, 287.7139, 287.7285, 287.7432, 287.7578, 
    287.7722, 287.7732, 287.7605, 287.7476, 287.7346, 287.7219, 287.709, 
    287.6963, 287.6833, 287.6707, 287.6577, 287.645, 287.6321, 287.6194, 
    287.5752, 287.5247, 287.4663, 287.3977, 287.3162, 287.2178, 287.0964, 
    286.9434, 285.2285, 285.1653, 285.1108, 285.0637, 284.9004, 284.6157, 
    284.3313, 284.0469, 283.7622, 283.4778, 283.1934, 282.9087, 282.6243, 
    282.3398, 282.0552, 281.7708, 281.4863, 281.511, 281.5356, 281.5605, 
    281.5852, 281.6099, 281.6348, 281.6594, 281.6841, 281.7087, 281.7336, 
    281.7583, 281.783, 281.7708, 281.7217, 281.6726, 281.6235, 281.5745, 
    281.5254, 281.4763, 281.4272, 281.3779, 281.3289, 281.2798, 281.2307, 
    281.1816, 281.1414, 281.1011, 281.0608, 281.0205, 280.9802, 280.9399, 
    280.8997, 280.8594, 280.8191, 280.7788, 280.7385, 280.6982, 280.666, 
    280.6423, 280.6184, 280.5945, 280.5708, 280.5469, 280.5229, 280.499, 
    280.4753, 280.4514, 280.4275, 280.4038, 280.3799, 280.3381, 280.2966, 
    280.2551, 280.2134, 280.1719, 280.1301, 280.0886, 280.0469, 280.0054, 
    279.9639, 279.9221, 279.8806, 279.8276, 279.7637, 279.6997, 279.6357, 
    279.5715, 279.5076, 279.4436, 279.3796, 279.3157, 279.2515, 279.1875, 
    279.1235, 279.0596, 279.0056, 278.9514, 278.8975, 278.8435, 278.7896, 
    278.7354, 278.6814, 278.6274, 278.5735, 278.5193, 278.4653, 278.4114, 
    278.3997, 278.4302, 278.4609, 278.4915, 278.522, 278.5525, 278.5833, 
    278.6138, 278.6443, 278.6748, 278.7056, 278.7361, 278.7666,
  287.0439, 287.1147, 287.1858, 287.2566, 287.3274, 287.3984, 287.4692, 
    287.54, 287.6111, 287.6819, 287.7527, 287.7961, 287.8396, 287.8831, 
    287.9268, 287.9702, 288.0137, 288.0571, 288.1006, 288.144, 288.1875, 
    288.231, 288.2744, 288.2993, 288.3052, 288.3113, 288.3174, 288.3235, 
    288.3296, 288.3357, 288.3416, 288.3477, 288.3538, 288.3599, 288.366, 
    288.3721, 288.3669, 288.3618, 288.3564, 288.3513, 288.3462, 288.3411, 
    288.3359, 288.3308, 288.3257, 288.3206, 288.3154, 288.3103, 288.3037, 
    288.2957, 288.2876, 288.2798, 288.2717, 288.2637, 288.2556, 288.2476, 
    288.2395, 288.2314, 288.2234, 288.2153, 288.2075, 288.2041, 288.2009, 
    288.1975, 288.1943, 288.1912, 288.1877, 288.1846, 288.1814, 288.178, 
    288.1748, 288.1716, 288.1682, 288.1416, 288.0918, 288.0417, 287.9917, 
    287.9419, 287.8918, 287.8418, 287.792, 287.7419, 287.6919, 287.6421, 
    287.592, 287.5422, 287.5261, 287.5103, 287.4941, 287.4783, 287.4624, 
    287.4463, 287.4304, 287.4146, 287.3984, 287.3826, 287.3667, 287.3506, 
    287.3442, 287.3474, 287.3503, 287.3535, 287.3567, 287.3596, 287.3628, 
    287.3657, 287.3689, 287.3721, 287.375, 287.3782, 287.3813, 287.3635, 
    287.3457, 287.3276, 287.3098, 287.292, 287.2742, 287.2563, 287.2385, 
    287.2207, 287.2029, 287.1851, 287.1672, 287.1768, 287.2141, 287.2512, 
    287.2886, 287.3257, 287.363, 287.4001, 287.4375, 287.4746, 287.512, 
    287.5491, 287.5864, 287.6235, 287.6379, 287.6521, 287.6665, 287.6807, 
    287.6948, 287.7092, 287.7234, 287.7378, 287.752, 287.7661, 287.7805, 
    287.7947, 287.7986, 287.7917, 287.7849, 287.7783, 287.7715, 287.7649, 
    287.7581, 287.7515, 287.7446, 287.7378, 287.7312, 287.7244, 287.7178, 
    287.6777, 287.6318, 287.5786, 287.5164, 287.4424, 287.353, 287.2427, 
    287.1038, 285.5459, 285.4885, 285.4392, 285.3965, 285.2197, 284.9053, 
    284.5908, 284.2764, 283.9619, 283.6475, 283.333, 283.0186, 282.7041, 
    282.3896, 282.0752, 281.7607, 281.4463, 281.47, 281.4934, 281.5171, 
    281.5408, 281.5645, 281.5879, 281.6116, 281.6353, 281.6589, 281.6824, 
    281.7061, 281.7297, 281.7178, 281.6702, 281.6228, 281.5752, 281.5278, 
    281.4805, 281.4329, 281.3855, 281.3379, 281.2905, 281.2429, 281.1956, 
    281.1479, 281.1082, 281.0684, 281.0283, 280.9885, 280.9485, 280.9087, 
    280.8689, 280.8289, 280.7891, 280.749, 280.7092, 280.6694, 280.6367, 
    280.6116, 280.5864, 280.5613, 280.5359, 280.5107, 280.4856, 280.4604, 
    280.4351, 280.4099, 280.3848, 280.3594, 280.3342, 280.2937, 280.2529, 
    280.2124, 280.1719, 280.1311, 280.0906, 280.0498, 280.0093, 279.9685, 
    279.928, 279.8875, 279.8467, 279.7952, 279.7329, 279.6707, 279.6082, 
    279.5459, 279.4836, 279.4211, 279.3589, 279.2966, 279.2344, 279.1719, 
    279.1096, 279.0474, 278.9946, 278.9419, 278.8892, 278.8364, 278.7837, 
    278.7312, 278.6785, 278.6257, 278.573, 278.5203, 278.4675, 278.4148, 
    278.3989, 278.4199, 278.4407, 278.4617, 278.4827, 278.5034, 278.5244, 
    278.5452, 278.5662, 278.5869, 278.6079, 278.6289, 278.6497 ;
}
